module top ( in0,  in1,  in2,  in3,  in4,  in5,  in6,  in7 , y1, y2 );

input in0,  in1,  in2,  in3, in4,  in5,  in6,  in7;
wire a , b , c , d, e, f;
output y1 , y2 ;
wire w1 , w2 , w3 , w4 , w5;
wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576;

nor ( n0, in0, in1 );
and ( n1, in0, in2 );
nor ( n2, in0, in3 );
xor ( n3, in0, in4 );
nor ( n4, in0, in5 );
and ( n5, in0, in6 );
nand ( n6, in0, in7 );
nand ( n7, in1, in2 );
nor ( n8, in1, in3 );
nor ( n9, in1, in4 );
and ( n10, in1, in5 );
or ( n11, in1, in6 );
or ( n12, in1, in7 );
and ( n13, in2, in3 );
nor ( n14, in2, in4 );
xor ( n15, in2, in5 );
nor ( n16, in2, in6 );
and ( n17, in2, in7 );
or ( n18, in3, in4 );
nand ( n19, in3, in5 );
and ( n20, in3, in6 );
nand ( n21, in3, in7 );
or ( n22, in4, in5 );
xor ( n23, in4, in6 );
xor ( n24, in4, in7 );
nand ( n25, in5, in6 );
xor ( n26, in5, in7 );
and ( n27, in6, in7 );
or ( n28, n6, n22 );
nand ( n29, n2, n16 );
xor ( n30, n4, n19 );
and ( n31, n5, n26 );
nor ( n32, n4, n13 );
and ( n33, n0, n8 );
or ( n34, n1, n21 );
nor ( n35, n15, n22 );
and ( n36, n1, n4 );
and ( n37, n5, n11 );
and ( n38, n19, n22 );
nand ( n39, n3, n24 );
or ( n40, n5, n12 );
and ( n41, n4, n15 );
nand ( n42, n2, n24 );
xor ( n43, n2, n22 );
or ( n44, n10, n17 );
nand ( n45, n13, n26 );
nor ( n46, n3, n7 );
nor ( n47, n9, n24 );
nor ( n48, n10, n11 );
or ( n49, n23, n24 );
and ( n50, n10, n24 );
xor ( n51, n9, n18 );
nand ( n52, n11, n23 );
xor ( n53, n7, n25 );
xor ( n54, n2, n26 );
xor ( n55, n8, n11 );
and ( n56, n10, n18 );
xor ( n57, n12, n19 );
and ( n58, n5, n20 );
nor ( n59, n21, n25 );
or ( n60, n0, n12 );
nor ( n61, n20, n21 );
or ( n62, n11, n18 );
nor ( n63, n4, n21 );
and ( n64, n1, n15 );
xor ( n65, n1, n12 );
or ( n66, n10, n20 );
and ( n67, n0, n25 );
or ( n68, n3, n18 );
xor ( n69, n10, n25 );
nand ( n70, n2, n4 );
nand ( n71, n11, n21 );
or ( n72, n2, n17 );
nand ( n73, n25, n26 );
nor ( n74, n11, n17 );
nor ( n75, n7, n13 );
or ( n76, n17, n22 );
or ( n77, n6, n20 );
nand ( n78, n2, n15 );
nand ( n79, n0, n6 );
xor ( n80, n16, n19 );
xor ( n81, n17, n19 );
xor ( n82, n6, n17 );
nand ( n83, n4, n12 );
xor ( n84, n4, n26 );
or ( n85, n7, n21 );
xor ( n86, n0, n17 );
nor ( n87, n18, n24 );
xor ( n88, n15, n25 );
nand ( n89, n9, n26 );
and ( n90, n11, n12 );
nor ( n91, n7, n24 );
or ( n92, n3, n9 );
xor ( n93, n0, n10 );
nand ( n94, n8, n13 );
or ( n95, n1, n8 );
xor ( n96, n9, n21 );
xor ( n97, n7, n17 );
and ( n98, n9, n19 );
nor ( n99, n9, n14 );
xor ( n100, n12, n26 );
nor ( n101, n18, n26 );
xor ( n102, n8, n19 );
nor ( n103, n14, n26 );
xor ( n104, n20, n26 );
and ( n105, n8, n25 );
or ( n106, n3, n5 );
and ( n107, n3, n22 );
and ( n108, n10, n14 );
nand ( n109, n4, n10 );
and ( n110, n11, n15 );
xor ( n111, n9, n11 );
nor ( n112, n3, n6 );
nor ( n113, n12, n17 );
nor ( n114, n2, n23 );
xor ( n115, n9, n13 );
nand ( n116, n12, n21 );
or ( n117, n6, n24 );
nand ( n118, n11, n13 );
and ( n119, n11, n19 );
xor ( n120, n14, n20 );
or ( n121, n11, n16 );
xor ( n122, n13, n18 );
and ( n123, n12, n18 );
or ( n124, n11, n25 );
nand ( n125, n8, n10 );
nand ( n126, n3, n12 );
nor ( n127, n4, n18 );
or ( n128, n5, n7 );
or ( n129, n21, n26 );
xor ( n130, n17, n25 );
nand ( n131, n18, n21 );
or ( n132, n2, n6 );
or ( n133, n8, n21 );
or ( n134, n6, n12 );
and ( n135, n3, n23 );
xor ( n136, n12, n20 );
nor ( n137, n2, n12 );
xor ( n138, n4, n17 );
xor ( n139, n22, n23 );
or ( n140, n4, n14 );
or ( n141, n1, n9 );
xor ( n142, n3, n19 );
nor ( n143, n2, n7 );
nand ( n144, n10, n13 );
or ( n145, n9, n17 );
and ( n146, n2, n57 );
or ( n147, n55, n86 );
nor ( n148, n126, n142 );
nor ( n149, n56, n96 );
nor ( n150, n42, n120 );
or ( n151, n14, n109 );
xor ( n152, n74, n125 );
or ( n153, n73, n97 );
xor ( n154, n5, n37 );
or ( n155, n29, n102 );
nor ( n156, n34, n89 );
xor ( n157, n23, n54 );
and ( n158, n77, n92 );
nand ( n159, n35, n80 );
nand ( n160, n4, n38 );
nor ( n161, n50, n132 );
and ( n162, n6, n89 );
nand ( n163, n7, n61 );
or ( n164, n5, n9 );
nand ( n165, n79, n89 );
xor ( n166, n37, n94 );
xor ( n167, n10, n137 );
xor ( n168, n49, n97 );
or ( n169, n14, n43 );
xor ( n170, n34, n53 );
xor ( n171, n70, n133 );
nand ( n172, n122, n127 );
nand ( n173, n49, n64 );
xor ( n174, n94, n111 );
nor ( n175, n10, n32 );
or ( n176, n105, n108 );
nor ( n177, n6, n92 );
or ( n178, n92, n104 );
xor ( n179, n81, n127 );
nor ( n180, n6, n72 );
xor ( n181, n44, n96 );
or ( n182, n44, n89 );
and ( n183, n89, n102 );
or ( n184, n120, n127 );
or ( n185, n78, n140 );
and ( n186, n49, n139 );
xor ( n187, n69, n92 );
nor ( n188, n29, n91 );
nor ( n189, n33, n53 );
nor ( n190, n19, n103 );
nor ( n191, n60, n108 );
or ( n192, n41, n127 );
or ( n193, n9, n42 );
or ( n194, n63, n97 );
nand ( n195, n3, n135 );
nand ( n196, n99, n143 );
or ( n197, n21, n109 );
xor ( n198, n69, n82 );
and ( n199, n62, n131 );
and ( n200, n9, n140 );
nor ( n201, n16, n78 );
and ( n202, n24, n103 );
nand ( n203, n7, n14 );
nand ( n204, n100, n113 );
nor ( n205, n42, n138 );
nor ( n206, n113, n139 );
and ( n207, n48, n113 );
and ( n208, n19, n130 );
nand ( n209, n73, n120 );
nand ( n210, n14, n132 );
and ( n211, n42, n96 );
nand ( n212, n2, n37 );
xor ( n213, n41, n64 );
xor ( n214, n67, n128 );
nand ( n215, n30, n107 );
or ( n216, n28, n118 );
xor ( n217, n88, n122 );
and ( n218, n2, n120 );
and ( n219, n58, n59 );
nand ( n220, n72, n108 );
or ( n221, n9, n86 );
nor ( n222, n3, n59 );
or ( n223, n61, n108 );
or ( n224, n45, n83 );
or ( n225, n14, n127 );
nor ( n226, n96, n107 );
or ( n227, n23, n25 );
xor ( n228, n54, n131 );
xor ( n229, n124, n130 );
nor ( n230, n63, n95 );
and ( n231, n69, n76 );
and ( n232, n6, n30 );
xor ( n233, n26, n109 );
nor ( n234, n11, n52 );
nor ( n235, n90, n138 );
nand ( n236, n2, n102 );
or ( n237, n3, n100 );
nor ( n238, n66, n135 );
and ( n239, n121, n122 );
xor ( n240, n16, n27 );
xor ( n241, n26, n57 );
nand ( n242, n2, n34 );
or ( n243, n60, n100 );
and ( n244, n81, n99 );
nor ( n245, n87, n139 );
xor ( n246, n2, n105 );
nor ( n247, n31, n89 );
or ( n248, n14, n100 );
xor ( n249, n32, n114 );
or ( n250, n12, n135 );
xor ( n251, n104, n142 );
and ( n252, n86, n132 );
and ( n253, n118, n135 );
nand ( n254, n25, n80 );
nand ( n255, n7, n40 );
nor ( n256, n132, n137 );
or ( n257, n14, n45 );
or ( n258, n29, n121 );
nor ( n259, n12, n126 );
and ( n260, n9, n95 );
xor ( n261, n94, n105 );
and ( n262, n32, n46 );
nor ( n263, n33, n129 );
and ( n264, n61, n90 );
nor ( n265, n65, n91 );
nand ( n266, n50, n131 );
or ( n267, n90, n132 );
or ( n268, n62, n136 );
and ( n269, n80, n88 );
nor ( n270, n63, n119 );
nand ( n271, n15, n143 );
or ( n272, n24, n50 );
nor ( n273, n1, n21 );
and ( n274, n1, n132 );
xor ( n275, n39, n107 );
nand ( n276, n50, n120 );
and ( n277, n25, n127 );
xor ( n278, n24, n72 );
nor ( n279, n107, n118 );
nor ( n280, n11, n73 );
xor ( n281, n7, n98 );
nand ( n282, n19, n128 );
nand ( n283, n61, n135 );
or ( n284, n1, n49 );
and ( n285, n71, n134 );
nand ( n286, n41, n90 );
xor ( n287, n73, n130 );
nand ( n288, n115, n125 );
or ( n289, n8, n35 );
xor ( n290, n71, n84 );
and ( n291, n24, n111 );
or ( n292, n73, n133 );
xor ( n293, n23, n93 );
nor ( n294, n70, n131 );
and ( n295, n43, n53 );
and ( n296, n18, n51 );
nand ( n297, n12, n141 );
nand ( n298, n20, n142 );
nor ( n299, n23, n37 );
xor ( n300, n8, n89 );
or ( n301, n74, n126 );
xor ( n302, n82, n105 );
and ( n303, n13, n42 );
nand ( n304, n2, n51 );
or ( n305, n57, n131 );
nand ( n306, n117, n122 );
or ( n307, n1, n18 );
nor ( n308, n87, n95 );
xor ( n309, n32, n45 );
xor ( n310, n56, n124 );
and ( n311, n71, n125 );
and ( n312, n81, n107 );
nand ( n313, n72, n121 );
nor ( n314, n70, n128 );
xor ( n315, n0, n19 );
and ( n316, n32, n44 );
nand ( n317, n27, n90 );
xor ( n318, n49, n82 );
xor ( n319, n47, n125 );
and ( n320, n58, n98 );
and ( n321, n40, n140 );
nor ( n322, n88, n96 );
and ( n323, n107, n132 );
or ( n324, n129, n133 );
or ( n325, n66, n132 );
and ( n326, n53, n82 );
or ( n327, n58, n107 );
nand ( n328, n51, n55 );
xor ( n329, n48, n88 );
nand ( n330, n20, n22 );
and ( n331, n23, n94 );
xor ( n332, n0, n132 );
nor ( n333, n59, n108 );
xor ( n334, n0, n61 );
or ( n335, n14, n37 );
or ( n336, n9, n38 );
nand ( n337, n65, n84 );
nand ( n338, n90, n100 );
and ( n339, n119, n126 );
and ( n340, n112, n140 );
and ( n341, n4, n78 );
or ( n342, n67, n136 );
and ( n343, n73, n91 );
nand ( n344, n74, n117 );
and ( n345, n4, n20 );
and ( n346, n18, n118 );
and ( n347, n42, n49 );
or ( n348, n23, n72 );
nor ( n349, n92, n132 );
or ( n350, n61, n122 );
xor ( n351, n3, n37 );
nand ( n352, n55, n66 );
xor ( n353, n111, n129 );
and ( n354, n100, n136 );
nor ( n355, n93, n102 );
and ( n356, n93, n133 );
xor ( n357, n49, n95 );
xor ( n358, n13, n129 );
and ( n359, n33, n89 );
nor ( n360, n10, n63 );
xor ( n361, n86, n95 );
and ( n362, n38, n73 );
nor ( n363, n18, n20 );
and ( n364, n55, n140 );
or ( n365, n25, n96 );
nor ( n366, n69, n81 );
nand ( n367, n112, n119 );
nor ( n368, n75, n79 );
nand ( n369, n34, n86 );
nor ( n370, n53, n63 );
xor ( n371, n1, n99 );
xor ( n372, n119, n130 );
or ( n373, n42, n109 );
and ( n374, n100, n122 );
and ( n375, n114, n138 );
and ( n376, n94, n122 );
or ( n377, n58, n139 );
and ( n378, n30, n66 );
nor ( n379, n7, n95 );
or ( n380, n39, n93 );
xor ( n381, n59, n138 );
or ( n382, n12, n88 );
and ( n383, n3, n39 );
nand ( n384, n54, n136 );
nor ( n385, n0, n42 );
or ( n386, n3, n43 );
and ( n387, n51, n62 );
nor ( n388, n59, n125 );
nand ( n389, n49, n132 );
or ( n390, n92, n95 );
nor ( n391, n99, n132 );
or ( n392, n27, n134 );
xor ( n393, n23, n119 );
nor ( n394, n75, n104 );
or ( n395, n62, n114 );
xor ( n396, n28, n128 );
nor ( n397, n6, n75 );
nand ( n398, n19, n91 );
or ( n399, n0, n104 );
xor ( n400, n69, n79 );
and ( n401, n59, n68 );
nor ( n402, n66, n118 );
nor ( n403, n89, n104 );
or ( n404, n37, n136 );
xor ( n405, n32, n40 );
xor ( n406, n52, n84 );
nand ( n407, n66, n86 );
nand ( n408, n106, n127 );
xor ( n409, n69, n102 );
or ( n410, n63, n106 );
or ( n411, n30, n123 );
nor ( n412, n44, n55 );
nor ( n413, n67, n114 );
nand ( n414, n99, n109 );
nor ( n415, n123, n125 );
xor ( n416, n17, n105 );
and ( n417, n7, n136 );
and ( n418, n53, n133 );
and ( n419, n52, n134 );
nand ( n420, n0, n11 );
nand ( n421, n70, n87 );
and ( n422, n20, n67 );
nor ( n423, n62, n79 );
nor ( n424, n2, n28 );
and ( n425, n56, n85 );
or ( n426, n13, n101 );
xor ( n427, n20, n31 );
or ( n428, n11, n94 );
xor ( n429, n41, n48 );
xor ( n430, n36, n37 );
nor ( n431, n51, n143 );
nor ( n432, n109, n111 );
and ( n433, n39, n139 );
and ( n434, n5, n40 );
xor ( n435, n80, n90 );
and ( n436, n117, n138 );
and ( n437, n7, n16 );
or ( n438, n83, n130 );
or ( n439, n128, n133 );
nor ( n440, n54, n71 );
and ( n441, n29, n46 );
nor ( n442, n103, n141 );
or ( n443, n50, n72 );
nor ( n444, n100, n138 );
xor ( n445, n66, n103 );
nor ( n446, n30, n31 );
xor ( n447, n63, n133 );
xor ( n448, n79, n143 );
nand ( n449, n96, n141 );
nand ( n450, n38, n65 );
nand ( n451, n8, n114 );
nor ( n452, n95, n117 );
xor ( n453, n42, n50 );
nor ( n454, n35, n125 );
nand ( n455, n68, n138 );
nor ( n456, n39, n57 );
or ( n457, n26, n95 );
nor ( n458, n39, n123 );
nor ( n459, n34, n61 );
nor ( n460, n25, n50 );
or ( n461, n80, n91 );
or ( n462, n95, n125 );
nor ( n463, n32, n107 );
nor ( n464, n18, n142 );
or ( n465, n55, n61 );
xor ( n466, n118, n136 );
xor ( n467, n25, n48 );
nor ( n468, n1, n121 );
nand ( n469, n80, n95 );
nor ( n470, n6, n87 );
nand ( n471, n28, n83 );
xor ( n472, n72, n130 );
and ( n473, n51, n108 );
nor ( n474, n67, n117 );
nor ( n475, n129, n136 );
xor ( n476, n77, n82 );
nand ( n477, n111, n118 );
or ( n478, n51, n99 );
or ( n479, n117, n121 );
xor ( n480, n58, n75 );
nand ( n481, n16, n60 );
or ( n482, n43, n90 );
and ( n483, n23, n74 );
xor ( n484, n25, n134 );
nand ( n485, n13, n79 );
nor ( n486, n6, n114 );
nor ( n487, n1, n134 );
and ( n488, n47, n139 );
or ( n489, n18, n23 );
or ( n490, n1, n69 );
and ( n491, n36, n142 );
nor ( n492, n50, n65 );
nand ( n493, n7, n118 );
xor ( n494, n6, n117 );
and ( n495, n114, n125 );
nand ( n496, n27, n115 );
nand ( n497, n14, n108 );
xor ( n498, n58, n78 );
nor ( n499, n38, n45 );
xor ( n500, n8, n44 );
nor ( n501, n118, n132 );
nor ( n502, n64, n93 );
nor ( n503, n8, n103 );
and ( n504, n17, n40 );
and ( n505, n55, n68 );
or ( n506, n44, n54 );
nand ( n507, n57, n103 );
nand ( n508, n83, n114 );
or ( n509, n20, n36 );
and ( n510, n41, n130 );
and ( n511, n98, n109 );
nand ( n512, n43, n111 );
and ( n513, n62, n140 );
xor ( n514, n52, n92 );
nor ( n515, n8, n36 );
nor ( n516, n91, n132 );
or ( n517, n52, n71 );
and ( n518, n53, n142 );
and ( n519, n15, n89 );
or ( n520, n102, n142 );
or ( n521, n29, n43 );
nor ( n522, n16, n34 );
nor ( n523, n0, n2 );
nand ( n524, n1, n6 );
nand ( n525, n34, n122 );
xor ( n526, n57, n80 );
or ( n527, n25, n94 );
or ( n528, n51, n130 );
nand ( n529, n46, n89 );
or ( n530, n20, n113 );
or ( n531, n62, n143 );
or ( n532, n69, n110 );
xor ( n533, n41, n116 );
or ( n534, n22, n93 );
nand ( n535, n114, n115 );
or ( n536, n52, n69 );
or ( n537, n46, n72 );
nand ( n538, n3, n18 );
or ( n539, n49, n71 );
nor ( n540, n26, n32 );
and ( n541, n39, n140 );
nor ( n542, n78, n116 );
and ( n543, n103, n113 );
or ( n544, n56, n70 );
or ( n545, n55, n93 );
nand ( n546, n39, n128 );
nand ( n547, n56, n134 );
nor ( n548, n78, n101 );
nand ( n549, n141, n143 );
nand ( n550, n45, n124 );
or ( n551, n33, n112 );
or ( n552, n18, n61 );
or ( n553, n19, n24 );
nor ( n554, n20, n92 );
or ( n555, n43, n75 );
xor ( n556, n31, n143 );
and ( n557, n73, n82 );
and ( n558, n20, n77 );
nor ( n559, n65, n98 );
xor ( n560, n80, n81 );
nor ( n561, n113, n135 );
or ( n562, n94, n138 );
xor ( n563, n23, n102 );
and ( n564, n2, n13 );
nand ( n565, n25, n27 );
nand ( n566, n85, n109 );
or ( n567, n2, n118 );
xor ( n568, n8, n119 );
and ( n569, n79, n107 );
and ( n570, n30, n105 );
nor ( n571, n32, n109 );
and ( n572, n53, n54 );
nand ( n573, n50, n98 );
nor ( n574, n82, n107 );
nor ( n575, n44, n100 );
and ( n576, n34, n73 );
nor ( n577, n30, n89 );
or ( n578, n120, n142 );
or ( n579, n95, n133 );
and ( n580, n31, n64 );
xor ( n581, n15, n96 );
and ( n582, n116, n121 );
and ( n583, n107, n140 );
and ( n584, n33, n71 );
or ( n585, n46, n90 );
nor ( n586, n17, n87 );
and ( n587, n2, n81 );
and ( n588, n79, n120 );
xor ( n589, n78, n93 );
nand ( n590, n24, n84 );
nor ( n591, n24, n125 );
xor ( n592, n16, n64 );
xor ( n593, n54, n100 );
and ( n594, n71, n120 );
or ( n595, n73, n108 );
and ( n596, n13, n115 );
and ( n597, n64, n123 );
or ( n598, n11, n131 );
or ( n599, n40, n121 );
and ( n600, n12, n81 );
nand ( n601, n42, n137 );
xor ( n602, n27, n106 );
or ( n603, n32, n34 );
and ( n604, n107, n136 );
xor ( n605, n75, n100 );
or ( n606, n22, n133 );
or ( n607, n27, n65 );
or ( n608, n108, n142 );
or ( n609, n54, n138 );
or ( n610, n40, n135 );
or ( n611, n70, n95 );
nor ( n612, n7, n41 );
or ( n613, n39, n118 );
xor ( n614, n104, n136 );
xor ( n615, n3, n53 );
nor ( n616, n4, n6 );
nor ( n617, n102, n129 );
nor ( n618, n2, n94 );
nor ( n619, n108, n129 );
xor ( n620, n53, n86 );
and ( n621, n45, n73 );
xor ( n622, n73, n79 );
nor ( n623, n6, n50 );
xor ( n624, n79, n133 );
or ( n625, n91, n138 );
and ( n626, n116, n127 );
nor ( n627, n30, n139 );
or ( n628, n82, n136 );
and ( n629, n26, n143 );
xor ( n630, n2, n17 );
or ( n631, n7, n53 );
or ( n632, n42, n61 );
and ( n633, n17, n102 );
xor ( n634, n59, n116 );
nand ( n635, n66, n93 );
and ( n636, n14, n92 );
and ( n637, n79, n100 );
nor ( n638, n11, n82 );
nand ( n639, n97, n126 );
nor ( n640, n115, n138 );
xor ( n641, n16, n131 );
nand ( n642, n29, n93 );
nor ( n643, n24, n63 );
or ( n644, n35, n68 );
and ( n645, n72, n123 );
and ( n646, n12, n124 );
or ( n647, n37, n90 );
and ( n648, n61, n139 );
nor ( n649, n78, n108 );
xor ( n650, n82, n142 );
and ( n651, n47, n116 );
and ( n652, n37, n88 );
nand ( n653, n126, n141 );
nand ( n654, n61, n64 );
nand ( n655, n23, n89 );
xor ( n656, n5, n123 );
or ( n657, n59, n74 );
nand ( n658, n23, n32 );
xor ( n659, n30, n40 );
or ( n660, n31, n81 );
nand ( n661, n5, n83 );
nor ( n662, n32, n64 );
nor ( n663, n108, n110 );
and ( n664, n29, n138 );
and ( n665, n18, n50 );
nor ( n666, n34, n78 );
nand ( n667, n22, n78 );
nor ( n668, n15, n16 );
xor ( n669, n34, n65 );
xor ( n670, n36, n53 );
nand ( n671, n15, n112 );
nor ( n672, n32, n39 );
and ( n673, n64, n129 );
xor ( n674, n30, n74 );
xor ( n675, n29, n85 );
and ( n676, n11, n119 );
xor ( n677, n50, n143 );
nand ( n678, n74, n132 );
nand ( n679, n3, n17 );
or ( n680, n44, n61 );
or ( n681, n68, n81 );
xor ( n682, n49, n110 );
nor ( n683, n10, n42 );
and ( n684, n62, n142 );
and ( n685, n94, n112 );
or ( n686, n37, n77 );
xor ( n687, n34, n129 );
nand ( n688, n31, n91 );
nor ( n689, n5, n84 );
nor ( n690, n109, n140 );
nand ( n691, n33, n58 );
nor ( n692, n53, n68 );
nand ( n693, n18, n21 );
nand ( n694, n43, n137 );
xor ( n695, n9, n94 );
xor ( n696, n10, n57 );
nor ( n697, n43, n97 );
nand ( n698, n9, n99 );
or ( n699, n4, n18 );
xor ( n700, n20, n55 );
and ( n701, n89, n135 );
or ( n702, n112, n127 );
or ( n703, n8, n24 );
xor ( n704, n59, n87 );
or ( n705, n24, n85 );
nand ( n706, n93, n140 );
nand ( n707, n39, n90 );
nor ( n708, n41, n83 );
nor ( n709, n30, n100 );
or ( n710, n33, n37 );
and ( n711, n71, n77 );
or ( n712, n65, n143 );
and ( n713, n1, n113 );
and ( n714, n120, n125 );
xor ( n715, n65, n106 );
or ( n716, n49, n70 );
nand ( n717, n28, n34 );
and ( n718, n61, n111 );
and ( n719, n105, n127 );
nand ( n720, n83, n136 );
or ( n721, n11, n140 );
and ( n722, n15, n138 );
nand ( n723, n97, n135 );
and ( n724, n78, n115 );
and ( n725, n19, n22 );
nor ( n726, n24, n95 );
and ( n727, n21, n112 );
or ( n728, n89, n92 );
xor ( n729, n43, n78 );
xor ( n730, n49, n55 );
nor ( n731, n28, n131 );
nand ( n732, n2, n103 );
or ( n733, n25, n54 );
or ( n734, n36, n119 );
nor ( n735, n34, n94 );
xor ( n736, n15, n77 );
nor ( n737, n8, n28 );
nor ( n738, n46, n63 );
nand ( n739, n51, n56 );
or ( n740, n69, n111 );
nand ( n741, n105, n137 );
nand ( n742, n60, n102 );
xor ( n743, n11, n114 );
or ( n744, n1, n136 );
xor ( n745, n65, n134 );
xor ( n746, n48, n110 );
nand ( n747, n30, n56 );
or ( n748, n26, n92 );
and ( n749, n24, n30 );
nand ( n750, n18, n112 );
nand ( n751, n136, n137 );
nand ( n752, n137, n141 );
and ( n753, n29, n39 );
xor ( n754, n115, n128 );
and ( n755, n47, n120 );
and ( n756, n34, n100 );
and ( n757, n86, n128 );
nor ( n758, n85, n92 );
or ( n759, n91, n119 );
nand ( n760, n21, n125 );
or ( n761, n96, n113 );
nor ( n762, n3, n19 );
or ( n763, n11, n84 );
xor ( n764, n3, n36 );
xor ( n765, n44, n87 );
and ( n766, n87, n103 );
xor ( n767, n36, n116 );
or ( n768, n60, n105 );
or ( n769, n76, n93 );
nand ( n770, n83, n102 );
xor ( n771, n51, n89 );
xor ( n772, n35, n89 );
xor ( n773, n115, n127 );
and ( n774, n117, n129 );
xor ( n775, n52, n97 );
nor ( n776, n19, n106 );
and ( n777, n15, n76 );
and ( n778, n78, n126 );
or ( n779, n79, n141 );
nor ( n780, n4, n70 );
and ( n781, n57, n110 );
xor ( n782, n17, n72 );
xor ( n783, n1, n38 );
nand ( n784, n29, n92 );
nand ( n785, n71, n100 );
and ( n786, n57, n99 );
and ( n787, n72, n124 );
xor ( n788, n34, n91 );
xor ( n789, n22, n143 );
xor ( n790, n9, n45 );
nor ( n791, n18, n119 );
nand ( n792, n15, n39 );
and ( n793, n12, n122 );
and ( n794, n65, n108 );
and ( n795, n49, n142 );
and ( n796, n14, n112 );
nor ( n797, n30, n117 );
and ( n798, n10, n109 );
nand ( n799, n66, n112 );
and ( n800, n24, n58 );
and ( n801, n39, n82 );
and ( n802, n45, n60 );
and ( n803, n36, n82 );
or ( n804, n41, n79 );
nor ( n805, n29, n133 );
or ( n806, n18, n113 );
or ( n807, n44, n71 );
nor ( n808, n106, n122 );
nor ( n809, n86, n91 );
or ( n810, n72, n138 );
or ( n811, n52, n101 );
and ( n812, n68, n83 );
xor ( n813, n101, n123 );
xor ( n814, n9, n75 );
nand ( n815, n20, n138 );
or ( n816, n100, n114 );
nor ( n817, n94, n131 );
xor ( n818, n76, n139 );
xor ( n819, n93, n143 );
nand ( n820, n28, n116 );
nor ( n821, n71, n121 );
or ( n822, n33, n130 );
nand ( n823, n61, n71 );
and ( n824, n13, n124 );
or ( n825, n4, n96 );
nand ( n826, n29, n38 );
nand ( n827, n26, n33 );
nor ( n828, n119, n122 );
xor ( n829, n10, n130 );
nor ( n830, n104, n114 );
nand ( n831, n106, n115 );
nor ( n832, n68, n119 );
or ( n833, n53, n94 );
nand ( n834, n17, n30 );
nand ( n835, n41, n60 );
nand ( n836, n26, n122 );
xor ( n837, n58, n89 );
and ( n838, n58, n76 );
nor ( n839, n54, n110 );
nand ( n840, n61, n82 );
and ( n841, n46, n59 );
nand ( n842, n81, n104 );
or ( n843, n55, n130 );
nor ( n844, n49, n118 );
nand ( n845, n70, n139 );
or ( n846, n1, n110 );
nand ( n847, n92, n97 );
xor ( n848, n15, n114 );
nor ( n849, n100, n124 );
or ( n850, n26, n44 );
nand ( n851, n44, n97 );
and ( n852, n22, n95 );
and ( n853, n24, n140 );
xor ( n854, n57, n60 );
nor ( n855, n43, n61 );
or ( n856, n78, n90 );
or ( n857, n84, n112 );
or ( n858, n80, n130 );
nor ( n859, n60, n89 );
and ( n860, n47, n109 );
xor ( n861, n17, n114 );
and ( n862, n34, n105 );
nor ( n863, n4, n92 );
nand ( n864, n39, n54 );
or ( n865, n50, n52 );
nor ( n866, n18, n143 );
nand ( n867, n50, n103 );
or ( n868, n7, n48 );
nand ( n869, n46, n49 );
or ( n870, n8, n98 );
xor ( n871, n9, n73 );
xor ( n872, n6, n66 );
nor ( n873, n91, n94 );
nand ( n874, n26, n130 );
or ( n875, n28, n82 );
and ( n876, n81, n138 );
nor ( n877, n108, n120 );
and ( n878, n74, n128 );
xor ( n879, n35, n44 );
nand ( n880, n52, n130 );
nor ( n881, n40, n84 );
and ( n882, n83, n105 );
nor ( n883, n6, n7 );
and ( n884, n14, n103 );
xor ( n885, n50, n124 );
xor ( n886, n45, n91 );
and ( n887, n25, n95 );
or ( n888, n63, n66 );
and ( n889, n29, n72 );
nor ( n890, n16, n49 );
or ( n891, n19, n100 );
xor ( n892, n35, n121 );
or ( n893, n25, n77 );
or ( n894, n2, n124 );
nand ( n895, n15, n40 );
xor ( n896, n11, n27 );
xor ( n897, n93, n109 );
nand ( n898, n3, n13 );
or ( n899, n81, n92 );
nand ( n900, n72, n107 );
xor ( n901, n68, n74 );
or ( n902, n3, n117 );
or ( n903, n10, n134 );
xor ( n904, n89, n91 );
and ( n905, n109, n141 );
nand ( n906, n36, n95 );
xor ( n907, n104, n127 );
and ( n908, n8, n91 );
xor ( n909, n17, n27 );
nor ( n910, n71, n80 );
and ( n911, n44, n103 );
or ( n912, n31, n131 );
xor ( n913, n26, n128 );
nand ( n914, n47, n66 );
and ( n915, n35, n115 );
xor ( n916, n3, n122 );
nand ( n917, n61, n106 );
xor ( n918, n35, n76 );
or ( n919, n57, n102 );
xor ( n920, n34, n133 );
nor ( n921, n85, n140 );
and ( n922, n29, n82 );
nor ( n923, n47, n55 );
and ( n924, n17, n126 );
or ( n925, n24, n65 );
and ( n926, n28, n76 );
or ( n927, n8, n20 );
or ( n928, n15, n53 );
xor ( n929, n15, n94 );
nand ( n930, n12, n65 );
xor ( n931, n110, n113 );
xor ( n932, n75, n94 );
nor ( n933, n61, n104 );
nor ( n934, n35, n98 );
and ( n935, n56, n75 );
xor ( n936, n51, n86 );
nor ( n937, n67, n112 );
and ( n938, n6, n126 );
or ( n939, n48, n70 );
nand ( n940, n5, n31 );
and ( n941, n25, n35 );
xor ( n942, n28, n130 );
nand ( n943, n17, n35 );
nor ( n944, n72, n140 );
nand ( n945, n83, n99 );
nand ( n946, n1, n62 );
xor ( n947, n70, n111 );
or ( n948, n60, n80 );
and ( n949, n85, n132 );
or ( n950, n47, n62 );
nand ( n951, n55, n91 );
and ( n952, n5, n59 );
or ( n953, n61, n94 );
nand ( n954, n36, n120 );
xor ( n955, n2, n14 );
and ( n956, n81, n94 );
or ( n957, n1, n124 );
or ( n958, n21, n22 );
nor ( n959, n98, n128 );
and ( n960, n3, n111 );
and ( n961, n108, n123 );
nor ( n962, n66, n71 );
xor ( n963, n66, n70 );
xor ( n964, n62, n115 );
and ( n965, n20, n114 );
xor ( n966, n8, n49 );
or ( n967, n38, n118 );
nor ( n968, n74, n106 );
or ( n969, n139, n140 );
nor ( n970, n117, n133 );
or ( n971, n43, n119 );
or ( n972, n53, n65 );
nor ( n973, n0, n1 );
nand ( n974, n60, n114 );
and ( n975, n62, n108 );
and ( n976, n77, n139 );
nor ( n977, n15, n142 );
or ( n978, n77, n106 );
xor ( n979, n86, n129 );
and ( n980, n120, n141 );
or ( n981, n38, n57 );
nor ( n982, n2, n3 );
xor ( n983, n73, n81 );
or ( n984, n14, n34 );
and ( n985, n47, n132 );
nand ( n986, n42, n70 );
nor ( n987, n45, n135 );
nor ( n988, n19, n137 );
xor ( n989, n56, n128 );
and ( n990, n17, n120 );
nand ( n991, n18, n136 );
nand ( n992, n67, n113 );
nor ( n993, n5, n36 );
and ( n994, n3, n68 );
nor ( n995, n54, n103 );
nor ( n996, n4, n110 );
or ( n997, n25, n108 );
and ( n998, n24, n98 );
and ( n999, n62, n96 );
nand ( n1000, n13, n93 );
or ( n1001, n137, n140 );
or ( n1002, n134, n142 );
xor ( n1003, n63, n118 );
nor ( n1004, n11, n55 );
nand ( n1005, n17, n138 );
nand ( n1006, n112, n138 );
and ( n1007, n44, n68 );
nor ( n1008, n6, n70 );
nand ( n1009, n14, n59 );
xor ( n1010, n76, n141 );
or ( n1011, n46, n127 );
nand ( n1012, n26, n41 );
or ( n1013, n26, n88 );
xor ( n1014, n57, n119 );
nor ( n1015, n117, n125 );
or ( n1016, n52, n117 );
xor ( n1017, n27, n39 );
and ( n1018, n26, n75 );
nor ( n1019, n12, n112 );
or ( n1020, n50, n91 );
and ( n1021, n13, n44 );
and ( n1022, n22, n115 );
and ( n1023, n56, n107 );
xor ( n1024, n40, n68 );
nor ( n1025, n53, n131 );
nor ( n1026, n17, n52 );
and ( n1027, n76, n87 );
nand ( n1028, n43, n74 );
or ( n1029, n12, n50 );
xor ( n1030, n14, n118 );
or ( n1031, n0, n47 );
xor ( n1032, n124, n131 );
or ( n1033, n62, n141 );
nand ( n1034, n120, n140 );
or ( n1035, n55, n138 );
nor ( n1036, n15, n119 );
or ( n1037, n97, n112 );
and ( n1038, n79, n86 );
nor ( n1039, n59, n65 );
and ( n1040, n63, n81 );
xor ( n1041, n117, n137 );
and ( n1042, n140, n143 );
xor ( n1043, n6, n12 );
xor ( n1044, n126, n136 );
xor ( n1045, n3, n32 );
nand ( n1046, n29, n40 );
and ( n1047, n19, n119 );
or ( n1048, n31, n58 );
and ( n1049, n8, n67 );
nand ( n1050, n97, n107 );
xor ( n1051, n3, n84 );
or ( n1052, n14, n89 );
xor ( n1053, n39, n122 );
xor ( n1054, n2, n143 );
or ( n1055, n8, n72 );
nor ( n1056, n85, n117 );
xor ( n1057, n71, n118 );
nand ( n1058, n49, n123 );
xor ( n1059, n50, n97 );
nor ( n1060, n3, n66 );
nor ( n1061, n30, n79 );
xor ( n1062, n50, n110 );
xor ( n1063, n1, n78 );
nand ( n1064, n94, n123 );
xor ( n1065, n43, n131 );
nand ( n1066, n11, n62 );
or ( n1067, n28, n68 );
xor ( n1068, n41, n53 );
nor ( n1069, n34, n127 );
and ( n1070, n0, n138 );
nor ( n1071, n113, n132 );
and ( n1072, n35, n46 );
and ( n1073, n5, n26 );
nand ( n1074, n55, n99 );
and ( n1075, n28, n132 );
xor ( n1076, n15, n128 );
xor ( n1077, n19, n127 );
or ( n1078, n49, n104 );
nand ( n1079, n40, n106 );
and ( n1080, n85, n126 );
or ( n1081, n37, n98 );
and ( n1082, n9, n114 );
or ( n1083, n64, n82 );
nand ( n1084, n57, n106 );
and ( n1085, n65, n105 );
nor ( n1086, n11, n89 );
nand ( n1087, n52, n100 );
nor ( n1088, n51, n82 );
nor ( n1089, n42, n112 );
xor ( n1090, n10, n126 );
nor ( n1091, n7, n15 );
and ( n1092, n128, n140 );
nor ( n1093, n118, n133 );
and ( n1094, n1, n116 );
and ( n1095, n34, n56 );
or ( n1096, n20, n71 );
and ( n1097, n28, n138 );
nor ( n1098, n14, n98 );
nor ( n1099, n42, n108 );
and ( n1100, n58, n108 );
nand ( n1101, n6, n24 );
nand ( n1102, n62, n124 );
xor ( n1103, n4, n129 );
nor ( n1104, n66, n85 );
nand ( n1105, n1, n70 );
nor ( n1106, n29, n119 );
nand ( n1107, n92, n133 );
or ( n1108, n61, n117 );
nand ( n1109, n79, n80 );
or ( n1110, n125, n136 );
nand ( n1111, n43, n46 );
nor ( n1112, n83, n115 );
nand ( n1113, n100, n102 );
xor ( n1114, n55, n136 );
nand ( n1115, n17, n81 );
nand ( n1116, n38, n58 );
nand ( n1117, n41, n56 );
nor ( n1118, n50, n56 );
nand ( n1119, n44, n116 );
or ( n1120, n75, n106 );
and ( n1121, n114, n139 );
nor ( n1122, n32, n41 );
nor ( n1123, n42, n88 );
and ( n1124, n88, n92 );
nor ( n1125, n45, n64 );
nand ( n1126, n81, n142 );
nand ( n1127, n18, n79 );
and ( n1128, n47, n110 );
nand ( n1129, n78, n91 );
xor ( n1130, n63, n109 );
xor ( n1131, n65, n104 );
xor ( n1132, n114, n130 );
nor ( n1133, n124, n126 );
nor ( n1134, n115, n123 );
and ( n1135, n6, n8 );
nor ( n1136, n18, n34 );
and ( n1137, n31, n45 );
and ( n1138, n33, n101 );
or ( n1139, n28, n105 );
nor ( n1140, n23, n80 );
or ( n1141, n3, n52 );
and ( n1142, n53, n137 );
xor ( n1143, n37, n44 );
xor ( n1144, n11, n57 );
xor ( n1145, n47, n122 );
nor ( n1146, n64, n105 );
xor ( n1147, n58, n136 );
xor ( n1148, n15, n90 );
xor ( n1149, n11, n24 );
and ( n1150, n1, n20 );
nor ( n1151, n59, n89 );
xor ( n1152, n41, n93 );
or ( n1153, n53, n119 );
nand ( n1154, n45, n109 );
and ( n1155, n45, n53 );
or ( n1156, n63, n125 );
and ( n1157, n113, n120 );
nand ( n1158, n94, n130 );
or ( n1159, n37, n99 );
nor ( n1160, n76, n86 );
xor ( n1161, n11, n50 );
nor ( n1162, n4, n17 );
nor ( n1163, n30, n90 );
or ( n1164, n20, n136 );
xor ( n1165, n14, n33 );
xor ( n1166, n102, n120 );
or ( n1167, n6, n84 );
nand ( n1168, n26, n116 );
xor ( n1169, n35, n116 );
or ( n1170, n44, n75 );
xor ( n1171, n110, n134 );
or ( n1172, n50, n142 );
and ( n1173, n23, n44 );
and ( n1174, n64, n100 );
or ( n1175, n78, n139 );
nand ( n1176, n4, n134 );
nor ( n1177, n78, n127 );
xor ( n1178, n80, n98 );
nand ( n1179, n122, n141 );
xor ( n1180, n46, n91 );
and ( n1181, n46, n93 );
or ( n1182, n60, n71 );
nand ( n1183, n12, n51 );
nand ( n1184, n80, n124 );
or ( n1185, n3, n15 );
xor ( n1186, n33, n95 );
or ( n1187, n18, n62 );
nor ( n1188, n3, n142 );
nor ( n1189, n51, n79 );
nand ( n1190, n61, n88 );
or ( n1191, n88, n115 );
xor ( n1192, n86, n130 );
nand ( n1193, n28, n57 );
nand ( n1194, n50, n140 );
xor ( n1195, n36, n41 );
nand ( n1196, n49, n79 );
or ( n1197, n65, n136 );
and ( n1198, n65, n119 );
nand ( n1199, n45, n119 );
and ( n1200, n108, n116 );
nor ( n1201, n19, n104 );
and ( n1202, n19, n69 );
or ( n1203, n20, n49 );
and ( n1204, n58, n106 );
nor ( n1205, n90, n118 );
nand ( n1206, n106, n125 );
or ( n1207, n78, n99 );
nor ( n1208, n92, n127 );
nand ( n1209, n59, n105 );
nor ( n1210, n56, n125 );
nor ( n1211, n37, n122 );
and ( n1212, n21, n111 );
nor ( n1213, n18, n116 );
and ( n1214, n48, n127 );
xor ( n1215, n9, n71 );
and ( n1216, n32, n35 );
nor ( n1217, n108, n118 );
or ( n1218, n53, n67 );
xor ( n1219, n21, n90 );
nor ( n1220, n40, n111 );
and ( n1221, n19, n134 );
nand ( n1222, n3, n89 );
or ( n1223, n85, n143 );
and ( n1224, n23, n90 );
nor ( n1225, n114, n122 );
and ( n1226, n24, n126 );
xor ( n1227, n8, n39 );
and ( n1228, n25, n115 );
and ( n1229, n59, n119 );
or ( n1230, n134, n139 );
nand ( n1231, n19, n73 );
and ( n1232, n31, n39 );
or ( n1233, n42, n83 );
xor ( n1234, n33, n92 );
or ( n1235, n33, n104 );
nor ( n1236, n31, n119 );
or ( n1237, n22, n77 );
nor ( n1238, n94, n135 );
nand ( n1239, n62, n139 );
or ( n1240, n88, n99 );
nand ( n1241, n17, n69 );
nor ( n1242, n107, n137 );
or ( n1243, n27, n95 );
or ( n1244, n9, n11 );
or ( n1245, n0, n60 );
or ( n1246, n98, n131 );
nor ( n1247, n93, n132 );
or ( n1248, n60, n140 );
nor ( n1249, n117, n130 );
xor ( n1250, n5, n89 );
nand ( n1251, n54, n117 );
or ( n1252, n33, n76 );
xor ( n1253, n122, n136 );
or ( n1254, n79, n98 );
xor ( n1255, n60, n88 );
nand ( n1256, n25, n65 );
nand ( n1257, n47, n95 );
nor ( n1258, n53, n56 );
and ( n1259, n73, n80 );
or ( n1260, n12, n86 );
nand ( n1261, n23, n103 );
and ( n1262, n13, n138 );
or ( n1263, n64, n92 );
and ( n1264, n35, n63 );
xor ( n1265, n0, n57 );
nand ( n1266, n57, n84 );
xor ( n1267, n14, n42 );
nor ( n1268, n5, n23 );
nor ( n1269, n5, n20 );
xor ( n1270, n63, n116 );
nor ( n1271, n7, n88 );
and ( n1272, n33, n61 );
nand ( n1273, n11, n51 );
or ( n1274, n37, n75 );
nand ( n1275, n29, n116 );
and ( n1276, n38, n81 );
nor ( n1277, n45, n127 );
nor ( n1278, n1, n25 );
nor ( n1279, n114, n116 );
xor ( n1280, n136, n140 );
or ( n1281, n47, n79 );
xor ( n1282, n59, n95 );
or ( n1283, n51, n83 );
or ( n1284, n44, n74 );
nand ( n1285, n16, n28 );
nand ( n1286, n39, n45 );
and ( n1287, n65, n116 );
and ( n1288, n16, n139 );
nand ( n1289, n17, n38 );
or ( n1290, n21, n115 );
nand ( n1291, n43, n135 );
or ( n1292, n3, n123 );
xor ( n1293, n59, n112 );
nand ( n1294, n55, n106 );
nor ( n1295, n46, n125 );
xor ( n1296, n4, n5 );
xor ( n1297, n47, n86 );
and ( n1298, n74, n97 );
and ( n1299, n0, n46 );
nor ( n1300, n79, n115 );
or ( n1301, n52, n67 );
or ( n1302, n78, n129 );
nand ( n1303, n92, n123 );
nand ( n1304, n43, n88 );
or ( n1305, n14, n86 );
xor ( n1306, n63, n89 );
nor ( n1307, n80, n96 );
nand ( n1308, n102, n131 );
xor ( n1309, n22, n82 );
and ( n1310, n32, n128 );
xor ( n1311, n12, n133 );
nor ( n1312, n66, n78 );
or ( n1313, n68, n72 );
nand ( n1314, n61, n138 );
or ( n1315, n27, n128 );
xor ( n1316, n91, n131 );
xor ( n1317, n58, n112 );
or ( n1318, n96, n119 );
nor ( n1319, n10, n121 );
nand ( n1320, n1, n91 );
or ( n1321, n20, n34 );
nand ( n1322, n39, n135 );
or ( n1323, n47, n72 );
or ( n1324, n89, n140 );
and ( n1325, n81, n115 );
xor ( n1326, n64, n111 );
nand ( n1327, n9, n100 );
and ( n1328, n5, n126 );
xor ( n1329, n81, n126 );
xor ( n1330, n89, n119 );
and ( n1331, n1, n87 );
and ( n1332, n34, n125 );
or ( n1333, n34, n119 );
xor ( n1334, n27, n141 );
nor ( n1335, n2, n58 );
and ( n1336, n71, n106 );
nor ( n1337, n16, n99 );
nor ( n1338, n38, n90 );
xor ( n1339, n124, n136 );
xor ( n1340, n98, n132 );
nor ( n1341, n32, n118 );
or ( n1342, n122, n134 );
xor ( n1343, n32, n141 );
and ( n1344, n10, n62 );
nand ( n1345, n31, n35 );
xor ( n1346, n57, n77 );
or ( n1347, n32, n36 );
xor ( n1348, n37, n95 );
nor ( n1349, n58, n82 );
xor ( n1350, n0, n117 );
nand ( n1351, n114, n137 );
or ( n1352, n40, n130 );
and ( n1353, n40, n81 );
xor ( n1354, n67, n106 );
and ( n1355, n11, n12 );
nor ( n1356, n110, n135 );
nor ( n1357, n17, n127 );
or ( n1358, n13, n70 );
and ( n1359, n0, n120 );
and ( n1360, n41, n115 );
nand ( n1361, n99, n138 );
or ( n1362, n4, n141 );
xor ( n1363, n19, n115 );
or ( n1364, n30, n54 );
nor ( n1365, n13, n131 );
and ( n1366, n7, n139 );
or ( n1367, n60, n94 );
xor ( n1368, n39, n87 );
nor ( n1369, n30, n49 );
or ( n1370, n5, n75 );
nor ( n1371, n71, n128 );
or ( n1372, n50, n102 );
or ( n1373, n129, n143 );
xor ( n1374, n4, n116 );
nand ( n1375, n61, n62 );
or ( n1376, n1, n31 );
xor ( n1377, n23, n95 );
nand ( n1378, n9, n28 );
xor ( n1379, n20, n86 );
xor ( n1380, n118, n128 );
and ( n1381, n5, n12 );
and ( n1382, n45, n54 );
xor ( n1383, n10, n26 );
nor ( n1384, n80, n114 );
or ( n1385, n19, n49 );
and ( n1386, n38, n76 );
xor ( n1387, n15, n95 );
nand ( n1388, n34, n132 );
xor ( n1389, n11, n121 );
nand ( n1390, n24, n31 );
nor ( n1391, n5, n139 );
xor ( n1392, n23, n107 );
and ( n1393, n57, n130 );
xor ( n1394, n15, n56 );
nor ( n1395, n18, n117 );
or ( n1396, n77, n118 );
nand ( n1397, n54, n96 );
nand ( n1398, n103, n134 );
nor ( n1399, n7, n52 );
or ( n1400, n15, n137 );
xor ( n1401, n65, n102 );
or ( n1402, n42, n52 );
nor ( n1403, n49, n135 );
and ( n1404, n72, n103 );
nand ( n1405, n47, n100 );
and ( n1406, n34, n70 );
or ( n1407, n23, n135 );
nor ( n1408, n68, n112 );
xor ( n1409, n31, n74 );
and ( n1410, n101, n135 );
xor ( n1411, n90, n127 );
xor ( n1412, n101, n121 );
or ( n1413, n47, n127 );
or ( n1414, n9, n112 );
and ( n1415, n8, n133 );
nand ( n1416, n22, n35 );
or ( n1417, n122, n139 );
nor ( n1418, n32, n70 );
and ( n1419, n36, n64 );
nand ( n1420, n18, n59 );
nand ( n1421, n35, n129 );
and ( n1422, n42, n51 );
and ( n1423, n0, n130 );
xor ( n1424, n37, n97 );
nor ( n1425, n24, n123 );
nor ( n1426, n75, n101 );
xor ( n1427, n24, n138 );
nand ( n1428, n51, n128 );
nand ( n1429, n45, n48 );
nor ( n1430, n101, n102 );
and ( n1431, n1, n139 );
nand ( n1432, n56, n66 );
or ( n1433, n94, n98 );
xor ( n1434, n119, n128 );
nor ( n1435, n49, n109 );
and ( n1436, n68, n141 );
nand ( n1437, n20, n62 );
or ( n1438, n58, n119 );
nand ( n1439, n117, n140 );
nor ( n1440, n8, n121 );
or ( n1441, n114, n119 );
and ( n1442, n41, n142 );
nor ( n1443, n25, n139 );
or ( n1444, n67, n129 );
nor ( n1445, n53, n83 );
nand ( n1446, n38, n119 );
nand ( n1447, n111, n142 );
or ( n1448, n39, n110 );
nor ( n1449, n85, n116 );
nand ( n1450, n14, n18 );
and ( n1451, n36, n141 );
or ( n1452, n13, n19 );
and ( n1453, n39, n46 );
and ( n1454, n105, n142 );
nand ( n1455, n33, n110 );
nor ( n1456, n19, n62 );
nand ( n1457, n7, n12 );
and ( n1458, n75, n142 );
or ( n1459, n16, n76 );
nor ( n1460, n4, n126 );
xor ( n1461, n10, n96 );
nor ( n1462, n56, n64 );
xor ( n1463, n13, n68 );
xor ( n1464, n31, n56 );
nor ( n1465, n75, n117 );
nand ( n1466, n46, n94 );
xor ( n1467, n38, n52 );
or ( n1468, n44, n48 );
nand ( n1469, n50, n119 );
or ( n1470, n20, n78 );
or ( n1471, n70, n74 );
nand ( n1472, n63, n88 );
xor ( n1473, n38, n139 );
and ( n1474, n89, n115 );
xor ( n1475, n5, n16 );
or ( n1476, n109, n129 );
nor ( n1477, n26, n63 );
or ( n1478, n77, n96 );
nand ( n1479, n56, n80 );
nand ( n1480, n10, n18 );
xor ( n1481, n22, n49 );
xor ( n1482, n77, n126 );
and ( n1483, n44, n124 );
xor ( n1484, n9, n91 );
xor ( n1485, n64, n118 );
nand ( n1486, n6, n60 );
and ( n1487, n60, n81 );
nand ( n1488, n102, n135 );
nand ( n1489, n24, n73 );
xor ( n1490, n9, n36 );
nand ( n1491, n124, n133 );
or ( n1492, n60, n74 );
or ( n1493, n84, n107 );
nand ( n1494, n79, n101 );
nand ( n1495, n91, n120 );
nor ( n1496, n54, n123 );
xor ( n1497, n57, n59 );
nor ( n1498, n116, n129 );
nand ( n1499, n43, n92 );
nand ( n1500, n100, n139 );
nor ( n1501, n79, n122 );
nor ( n1502, n107, n141 );
nand ( n1503, n88, n105 );
nand ( n1504, n35, n77 );
nor ( n1505, n60, n134 );
nand ( n1506, n130, n143 );
xor ( n1507, n50, n96 );
nor ( n1508, n82, n120 );
nor ( n1509, n78, n138 );
nand ( n1510, n66, n109 );
nor ( n1511, n113, n124 );
xor ( n1512, n43, n79 );
or ( n1513, n109, n120 );
xor ( n1514, n62, n88 );
and ( n1515, n74, n136 );
nor ( n1516, n28, n32 );
nand ( n1517, n82, n124 );
and ( n1518, n55, n101 );
xor ( n1519, n88, n117 );
xor ( n1520, n11, n32 );
and ( n1521, n37, n85 );
and ( n1522, n25, n140 );
nor ( n1523, n24, n139 );
nand ( n1524, n22, n111 );
or ( n1525, n58, n84 );
nor ( n1526, n102, n103 );
nor ( n1527, n36, n85 );
nor ( n1528, n0, n18 );
nor ( n1529, n5, n122 );
nor ( n1530, n51, n98 );
xor ( n1531, n67, n98 );
and ( n1532, n25, n107 );
nand ( n1533, n97, n104 );
or ( n1534, n37, n63 );
nand ( n1535, n128, n136 );
nor ( n1536, n55, n115 );
and ( n1537, n21, n84 );
or ( n1538, n45, n81 );
or ( n1539, n71, n117 );
nand ( n1540, n101, n131 );
and ( n1541, n46, n110 );
xor ( n1542, n23, n58 );
nand ( n1543, n18, n107 );
nand ( n1544, n5, n127 );
nor ( n1545, n127, n135 );
nand ( n1546, n21, n135 );
nor ( n1547, n56, n60 );
nor ( n1548, n34, n140 );
nor ( n1549, n60, n135 );
nor ( n1550, n2, n53 );
xor ( n1551, n27, n132 );
xor ( n1552, n43, n69 );
or ( n1553, n28, n137 );
nand ( n1554, n12, n128 );
nor ( n1555, n58, n92 );
nand ( n1556, n3, n41 );
xor ( n1557, n65, n80 );
or ( n1558, n25, n110 );
nand ( n1559, n2, n21 );
nor ( n1560, n57, n86 );
nand ( n1561, n113, n141 );
xor ( n1562, n120, n133 );
nand ( n1563, n53, n61 );
xor ( n1564, n26, n29 );
xor ( n1565, n44, n142 );
nand ( n1566, n101, n125 );
xor ( n1567, n123, n142 );
nor ( n1568, n76, n121 );
and ( n1569, n20, n43 );
nor ( n1570, n68, n128 );
nor ( n1571, n66, n94 );
xor ( n1572, n74, n120 );
xor ( n1573, n25, n136 );
xor ( n1574, n17, n82 );
nand ( n1575, n55, n121 );
xor ( n1576, n45, n61 );
nand ( n1577, n11, n122 );
and ( n1578, n12, n33 );
nand ( n1579, n7, n64 );
and ( n1580, n2, n20 );
nor ( n1581, n86, n115 );
or ( n1582, n62, n100 );
nor ( n1583, n66, n80 );
nand ( n1584, n113, n143 );
nand ( n1585, n28, n142 );
and ( n1586, n48, n101 );
and ( n1587, n64, n72 );
xor ( n1588, n11, n38 );
or ( n1589, n124, n139 );
nor ( n1590, n37, n113 );
and ( n1591, n4, n77 );
nor ( n1592, n53, n114 );
xor ( n1593, n31, n118 );
nand ( n1594, n27, n40 );
and ( n1595, n6, n37 );
xor ( n1596, n9, n35 );
and ( n1597, n45, n96 );
nand ( n1598, n57, n78 );
nor ( n1599, n64, n81 );
nor ( n1600, n20, n132 );
or ( n1601, n64, n87 );
and ( n1602, n8, n95 );
and ( n1603, n74, n134 );
nor ( n1604, n7, n101 );
nor ( n1605, n34, n120 );
or ( n1606, n75, n125 );
nand ( n1607, n65, n95 );
nor ( n1608, n54, n97 );
or ( n1609, n55, n134 );
nor ( n1610, n17, n93 );
xor ( n1611, n69, n119 );
nand ( n1612, n41, n51 );
xor ( n1613, n93, n138 );
nand ( n1614, n25, n87 );
nand ( n1615, n51, n87 );
and ( n1616, n80, n89 );
and ( n1617, n58, n86 );
or ( n1618, n112, n120 );
xor ( n1619, n36, n106 );
xor ( n1620, n30, n39 );
and ( n1621, n0, n44 );
or ( n1622, n2, n84 );
xor ( n1623, n88, n94 );
or ( n1624, n17, n78 );
nand ( n1625, n55, n94 );
xor ( n1626, n24, n40 );
nand ( n1627, n21, n72 );
nor ( n1628, n64, n114 );
xor ( n1629, n36, n136 );
or ( n1630, n40, n54 );
nand ( n1631, n11, n117 );
and ( n1632, n35, n43 );
and ( n1633, n2, n100 );
nand ( n1634, n22, n141 );
nor ( n1635, n44, n81 );
or ( n1636, n5, n118 );
nor ( n1637, n79, n95 );
or ( n1638, n1, n42 );
and ( n1639, n41, n73 );
nor ( n1640, n19, n45 );
xor ( n1641, n29, n106 );
xor ( n1642, n23, n143 );
nor ( n1643, n96, n108 );
xor ( n1644, n66, n141 );
nor ( n1645, n43, n60 );
or ( n1646, n56, n122 );
nand ( n1647, n3, n6 );
and ( n1648, n47, n104 );
nand ( n1649, n17, n65 );
nand ( n1650, n21, n141 );
and ( n1651, n72, n127 );
xor ( n1652, n75, n99 );
and ( n1653, n36, n115 );
nand ( n1654, n100, n117 );
and ( n1655, n96, n112 );
nor ( n1656, n33, n98 );
or ( n1657, n31, n53 );
nor ( n1658, n20, n56 );
nor ( n1659, n31, n84 );
or ( n1660, n112, n121 );
nor ( n1661, n22, n142 );
or ( n1662, n49, n106 );
or ( n1663, n60, n118 );
and ( n1664, n96, n140 );
and ( n1665, n9, n65 );
xor ( n1666, n24, n121 );
or ( n1667, n130, n131 );
nand ( n1668, n114, n123 );
nor ( n1669, n83, n129 );
xor ( n1670, n70, n81 );
or ( n1671, n9, n136 );
nor ( n1672, n1, n29 );
nand ( n1673, n31, n90 );
nand ( n1674, n57, n118 );
xor ( n1675, n91, n135 );
xor ( n1676, n32, n137 );
and ( n1677, n5, n66 );
or ( n1678, n94, n101 );
and ( n1679, n113, n138 );
nor ( n1680, n32, n63 );
xor ( n1681, n50, n54 );
xor ( n1682, n58, n87 );
and ( n1683, n30, n38 );
and ( n1684, n22, n97 );
xor ( n1685, n3, n101 );
or ( n1686, n23, n78 );
nor ( n1687, n21, n102 );
nand ( n1688, n31, n70 );
xor ( n1689, n40, n59 );
nand ( n1690, n28, n72 );
xor ( n1691, n80, n103 );
nand ( n1692, n24, n112 );
or ( n1693, n65, n123 );
and ( n1694, n43, n125 );
or ( n1695, n96, n98 );
nand ( n1696, n10, n112 );
nor ( n1697, n9, n18 );
nand ( n1698, n40, n134 );
nor ( n1699, n6, n48 );
and ( n1700, n43, n94 );
or ( n1701, n48, n69 );
xor ( n1702, n41, n72 );
and ( n1703, n23, n81 );
nand ( n1704, n11, n137 );
nand ( n1705, n58, n88 );
nand ( n1706, n27, n62 );
nand ( n1707, n22, n96 );
nand ( n1708, n55, n90 );
nand ( n1709, n44, n133 );
or ( n1710, n39, n92 );
xor ( n1711, n7, n99 );
and ( n1712, n28, n59 );
nand ( n1713, n35, n137 );
nor ( n1714, n23, n111 );
xor ( n1715, n69, n115 );
xor ( n1716, n68, n137 );
nor ( n1717, n7, n140 );
nand ( n1718, n16, n29 );
nor ( n1719, n26, n87 );
nor ( n1720, n26, n127 );
nor ( n1721, n6, n56 );
xor ( n1722, n74, n87 );
xor ( n1723, n61, n102 );
xor ( n1724, n24, n71 );
nor ( n1725, n49, n63 );
and ( n1726, n21, n94 );
nor ( n1727, n4, n125 );
xor ( n1728, n25, n109 );
or ( n1729, n8, n27 );
xor ( n1730, n1, n142 );
and ( n1731, n87, n90 );
and ( n1732, n113, n114 );
and ( n1733, n56, n67 );
and ( n1734, n17, n23 );
xor ( n1735, n0, n103 );
nand ( n1736, n86, n118 );
nand ( n1737, n71, n79 );
xor ( n1738, n97, n125 );
or ( n1739, n38, n122 );
xor ( n1740, n69, n133 );
or ( n1741, n136, n142 );
or ( n1742, n14, n101 );
nand ( n1743, n134, n140 );
nand ( n1744, n71, n90 );
nand ( n1745, n37, n114 );
nand ( n1746, n34, n43 );
and ( n1747, n38, n107 );
xor ( n1748, n58, n96 );
and ( n1749, n95, n103 );
nand ( n1750, n79, n85 );
and ( n1751, n14, n138 );
xor ( n1752, n132, n139 );
and ( n1753, n51, n53 );
nand ( n1754, n72, n129 );
and ( n1755, n73, n131 );
xor ( n1756, n1, n76 );
xor ( n1757, n46, n66 );
or ( n1758, n91, n126 );
or ( n1759, n27, n80 );
xor ( n1760, n69, n124 );
nand ( n1761, n69, n98 );
xor ( n1762, n90, n96 );
or ( n1763, n41, n88 );
and ( n1764, n1, n34 );
or ( n1765, n92, n136 );
nor ( n1766, n51, n136 );
nor ( n1767, n103, n136 );
nor ( n1768, n126, n137 );
nand ( n1769, n20, n108 );
nand ( n1770, n136, n138 );
and ( n1771, n82, n113 );
or ( n1772, n101, n107 );
nor ( n1773, n77, n137 );
and ( n1774, n48, n68 );
or ( n1775, n90, n101 );
nand ( n1776, n49, n66 );
xor ( n1777, n4, n119 );
nor ( n1778, n25, n41 );
or ( n1779, n79, n128 );
and ( n1780, n11, n47 );
or ( n1781, n15, n33 );
or ( n1782, n27, n51 );
xor ( n1783, n110, n129 );
and ( n1784, n47, n81 );
nand ( n1785, n0, n30 );
nor ( n1786, n90, n133 );
nand ( n1787, n90, n110 );
nor ( n1788, n119, n127 );
nor ( n1789, n14, n136 );
nand ( n1790, n15, n121 );
and ( n1791, n28, n45 );
or ( n1792, n119, n136 );
or ( n1793, n62, n92 );
or ( n1794, n41, n67 );
or ( n1795, n0, n112 );
nand ( n1796, n70, n135 );
and ( n1797, n29, n84 );
nand ( n1798, n83, n117 );
nor ( n1799, n8, n118 );
nand ( n1800, n54, n140 );
and ( n1801, n35, n133 );
nor ( n1802, n30, n112 );
and ( n1803, n17, n112 );
xor ( n1804, n22, n23 );
and ( n1805, n22, n92 );
and ( n1806, n36, n57 );
and ( n1807, n30, n68 );
and ( n1808, n43, n95 );
and ( n1809, n34, n87 );
xor ( n1810, n40, n102 );
or ( n1811, n86, n133 );
xor ( n1812, n82, n131 );
xor ( n1813, n5, n21 );
nor ( n1814, n41, n106 );
and ( n1815, n6, n55 );
nand ( n1816, n91, n121 );
or ( n1817, n73, n96 );
or ( n1818, n74, n105 );
and ( n1819, n3, n87 );
and ( n1820, n63, n93 );
or ( n1821, n8, n134 );
nand ( n1822, n9, n60 );
xor ( n1823, n57, n92 );
nor ( n1824, n19, n52 );
or ( n1825, n101, n128 );
or ( n1826, n125, n128 );
xor ( n1827, n89, n112 );
nand ( n1828, n39, n44 );
xor ( n1829, n62, n128 );
nor ( n1830, n114, n129 );
or ( n1831, n112, n136 );
nand ( n1832, n130, n141 );
nor ( n1833, n22, n138 );
nor ( n1834, n45, n74 );
nor ( n1835, n38, n68 );
or ( n1836, n42, n134 );
or ( n1837, n73, n87 );
xor ( n1838, n53, n87 );
or ( n1839, n8, n106 );
nor ( n1840, n13, n114 );
and ( n1841, n104, n125 );
or ( n1842, n63, n65 );
or ( n1843, n36, n137 );
nor ( n1844, n27, n129 );
or ( n1845, n33, n36 );
and ( n1846, n30, n60 );
and ( n1847, n49, n131 );
and ( n1848, n3, n44 );
and ( n1849, n5, n42 );
nand ( n1850, n10, n59 );
nor ( n1851, n12, n98 );
nand ( n1852, n22, n71 );
nor ( n1853, n105, n106 );
or ( n1854, n45, n56 );
nand ( n1855, n24, n53 );
nand ( n1856, n12, n28 );
nor ( n1857, n55, n95 );
nor ( n1858, n9, n26 );
or ( n1859, n27, n138 );
nor ( n1860, n28, n37 );
nor ( n1861, n18, n19 );
or ( n1862, n39, n72 );
or ( n1863, n27, n113 );
nor ( n1864, n23, n123 );
xor ( n1865, n67, n100 );
nor ( n1866, n108, n134 );
nand ( n1867, n99, n140 );
nand ( n1868, n22, n60 );
nor ( n1869, n6, n71 );
or ( n1870, n14, n125 );
and ( n1871, n96, n131 );
or ( n1872, n49, n127 );
nand ( n1873, n76, n117 );
or ( n1874, n82, n126 );
and ( n1875, n54, n141 );
nor ( n1876, n91, n127 );
and ( n1877, n129, n142 );
and ( n1878, n45, n105 );
and ( n1879, n59, n91 );
nand ( n1880, n106, n135 );
or ( n1881, n18, n132 );
nand ( n1882, n50, n100 );
or ( n1883, n7, n133 );
or ( n1884, n84, n97 );
xor ( n1885, n53, n66 );
and ( n1886, n15, n27 );
nor ( n1887, n76, n122 );
nor ( n1888, n16, n39 );
xor ( n1889, n35, n138 );
and ( n1890, n6, n90 );
xor ( n1891, n10, n11 );
xor ( n1892, n5, n72 );
nor ( n1893, n39, n96 );
nor ( n1894, n77, n100 );
nand ( n1895, n37, n82 );
and ( n1896, n79, n135 );
nor ( n1897, n12, n17 );
nor ( n1898, n98, n111 );
nand ( n1899, n21, n114 );
xor ( n1900, n108, n124 );
nand ( n1901, n75, n143 );
and ( n1902, n4, n109 );
and ( n1903, n7, n137 );
or ( n1904, n35, n60 );
nand ( n1905, n50, n55 );
xor ( n1906, n11, n85 );
nand ( n1907, n12, n27 );
nor ( n1908, n43, n142 );
or ( n1909, n2, n89 );
xor ( n1910, n7, n107 );
nand ( n1911, n59, n123 );
and ( n1912, n110, n117 );
or ( n1913, n81, n117 );
and ( n1914, n40, n47 );
nand ( n1915, n27, n79 );
nand ( n1916, n115, n131 );
and ( n1917, n114, n142 );
nor ( n1918, n8, n115 );
or ( n1919, n46, n61 );
nor ( n1920, n91, n125 );
nand ( n1921, n122, n140 );
and ( n1922, n0, n122 );
or ( n1923, n40, n131 );
nor ( n1924, n27, n78 );
nand ( n1925, n92, n142 );
nand ( n1926, n5, n138 );
xor ( n1927, n69, n78 );
nand ( n1928, n84, n121 );
nor ( n1929, n92, n130 );
xor ( n1930, n12, n123 );
xor ( n1931, n39, n40 );
xor ( n1932, n71, n129 );
nand ( n1933, n142, n143 );
nor ( n1934, n49, n73 );
or ( n1935, n102, n139 );
xor ( n1936, n111, n138 );
xor ( n1937, n12, n63 );
nor ( n1938, n108, n127 );
nor ( n1939, n33, n73 );
nand ( n1940, n18, n52 );
nor ( n1941, n40, n101 );
nor ( n1942, n31, n101 );
nand ( n1943, n29, n130 );
and ( n1944, n46, n70 );
or ( n1945, n0, n129 );
nand ( n1946, n3, n51 );
nand ( n1947, n90, n136 );
nand ( n1948, n105, n113 );
or ( n1949, n124, n135 );
nor ( n1950, n48, n125 );
nor ( n1951, n60, n129 );
nand ( n1952, n88, n141 );
xor ( n1953, n33, n59 );
nand ( n1954, n13, n110 );
xor ( n1955, n46, n113 );
nand ( n1956, n2, n131 );
nor ( n1957, n90, n131 );
nand ( n1958, n43, n84 );
and ( n1959, n24, n69 );
or ( n1960, n19, n32 );
or ( n1961, n98, n103 );
and ( n1962, n26, n100 );
nand ( n1963, n3, n125 );
nor ( n1964, n7, n66 );
nand ( n1965, n37, n93 );
and ( n1966, n7, n50 );
nor ( n1967, n75, n85 );
or ( n1968, n15, n26 );
xor ( n1969, n57, n121 );
or ( n1970, n85, n96 );
nor ( n1971, n99, n123 );
nand ( n1972, n80, n122 );
xor ( n1973, n2, n8 );
and ( n1974, n29, n110 );
or ( n1975, n1, n90 );
nor ( n1976, n43, n66 );
nor ( n1977, n72, n86 );
nand ( n1978, n9, n79 );
nor ( n1979, n59, n71 );
and ( n1980, n79, n126 );
and ( n1981, n69, n109 );
and ( n1982, n31, n141 );
xor ( n1983, n9, n23 );
and ( n1984, n29, n44 );
or ( n1985, n3, n14 );
nor ( n1986, n43, n108 );
nor ( n1987, n66, n102 );
nor ( n1988, n24, n137 );
nor ( n1989, n13, n82 );
or ( n1990, n19, n36 );
xor ( n1991, n1, n44 );
or ( n1992, n32, n47 );
or ( n1993, n111, n117 );
and ( n1994, n4, n83 );
nand ( n1995, n101, n108 );
xor ( n1996, n93, n112 );
and ( n1997, n135, n142 );
xor ( n1998, n35, n105 );
and ( n1999, n51, n80 );
and ( n2000, n91, n111 );
and ( n2001, n139, n143 );
nor ( n2002, n7, n59 );
nor ( n2003, n103, n118 );
xor ( n2004, n43, n83 );
and ( n2005, n56, n131 );
nor ( n2006, n36, n46 );
or ( n2007, n15, n59 );
nor ( n2008, n6, n125 );
nand ( n2009, n54, n119 );
and ( n2010, n21, n89 );
nor ( n2011, n72, n94 );
or ( n2012, n111, n122 );
nand ( n2013, n9, n87 );
xor ( n2014, n4, n34 );
xor ( n2015, n80, n140 );
and ( n2016, n78, n142 );
and ( n2017, n10, n66 );
and ( n2018, n35, n61 );
xor ( n2019, n38, n143 );
nand ( n2020, n67, n123 );
xor ( n2021, n8, n102 );
nand ( n2022, n8, n34 );
xor ( n2023, n111, n120 );
nor ( n2024, n40, n44 );
or ( n2025, n116, n131 );
xor ( n2026, n13, n116 );
xor ( n2027, n7, n111 );
nand ( n2028, n17, n89 );
or ( n2029, n113, n126 );
nand ( n2030, n113, n117 );
nand ( n2031, n75, n88 );
or ( n2032, n23, n99 );
nand ( n2033, n40, n126 );
nand ( n2034, n64, n78 );
or ( n2035, n33, n123 );
xor ( n2036, n55, n127 );
nor ( n2037, n116, n118 );
nor ( n2038, n88, n140 );
nor ( n2039, n101, n136 );
nor ( n2040, n50, n82 );
and ( n2041, n39, n100 );
nand ( n2042, n16, n19 );
xor ( n2043, n66, n131 );
nor ( n2044, n59, n113 );
and ( n2045, n38, n128 );
nand ( n2046, n57, n143 );
xor ( n2047, n23, n110 );
nor ( n2048, n75, n115 );
xor ( n2049, n17, n132 );
and ( n2050, n35, n56 );
or ( n2051, n66, n83 );
xor ( n2052, n47, n121 );
or ( n2053, n49, n83 );
xor ( n2054, n13, n122 );
nor ( n2055, n124, n127 );
or ( n2056, n2, n24 );
nor ( n2057, n0, n55 );
and ( n2058, n83, n119 );
or ( n2059, n36, n117 );
nor ( n2060, n77, n113 );
nand ( n2061, n25, n121 );
or ( n2062, n28, n86 );
xor ( n2063, n6, n31 );
nor ( n2064, n75, n112 );
xor ( n2065, n77, n119 );
nor ( n2066, n42, n75 );
nor ( n2067, n66, n67 );
nor ( n2068, n33, n52 );
and ( n2069, n75, n77 );
nand ( n2070, n37, n42 );
xor ( n2071, n47, n142 );
or ( n2072, n3, n30 );
nor ( n2073, n27, n118 );
nand ( n2074, n83, n94 );
nor ( n2075, n123, n133 );
nor ( n2076, n89, n111 );
nand ( n2077, n32, n91 );
and ( n2078, n14, n30 );
or ( n2079, n20, n124 );
nand ( n2080, n17, n106 );
nor ( n2081, n27, n84 );
or ( n2082, n40, n52 );
xor ( n2083, n13, n95 );
nor ( n2084, n62, n70 );
nor ( n2085, n10, n119 );
and ( n2086, n43, n117 );
nor ( n2087, n20, n74 );
and ( n2088, n5, n140 );
xor ( n2089, n47, n48 );
and ( n2090, n18, n26 );
nor ( n2091, n53, n89 );
nand ( n2092, n7, n81 );
nor ( n2093, n22, n125 );
nand ( n2094, n87, n91 );
or ( n2095, n31, n94 );
or ( n2096, n133, n139 );
nand ( n2097, n63, n121 );
or ( n2098, n18, n29 );
or ( n2099, n38, n74 );
and ( n2100, n20, n83 );
and ( n2101, n17, n45 );
nor ( n2102, n25, n38 );
nor ( n2103, n41, n133 );
xor ( n2104, n23, n39 );
xor ( n2105, n10, n13 );
xor ( n2106, n87, n97 );
or ( n2107, n65, n75 );
and ( n2108, n31, n125 );
nand ( n2109, n88, n128 );
xor ( n2110, n62, n93 );
nand ( n2111, n32, n50 );
xor ( n2112, n68, n133 );
or ( n2113, n4, n42 );
nand ( n2114, n40, n87 );
and ( n2115, n38, n66 );
nor ( n2116, n34, n41 );
xor ( n2117, n46, n108 );
or ( n2118, n53, n81 );
nor ( n2119, n28, n70 );
xor ( n2120, n27, n82 );
nor ( n2121, n97, n121 );
nor ( n2122, n22, n62 );
and ( n2123, n79, n84 );
xor ( n2124, n25, n76 );
nor ( n2125, n32, n53 );
nand ( n2126, n75, n118 );
xor ( n2127, n108, n109 );
and ( n2128, n23, n47 );
nand ( n2129, n5, n6 );
and ( n2130, n50, n134 );
nand ( n2131, n44, n114 );
xor ( n2132, n0, n96 );
and ( n2133, n3, n4 );
nand ( n2134, n19, n133 );
nand ( n2135, n12, n92 );
and ( n2136, n116, n135 );
xor ( n2137, n18, n104 );
nor ( n2138, n34, n77 );
nand ( n2139, n60, n104 );
nand ( n2140, n90, n103 );
nor ( n2141, n30, n138 );
xor ( n2142, n8, n63 );
nor ( n2143, n108, n140 );
and ( n2144, n55, n85 );
and ( n2145, n18, n65 );
and ( n2146, n58, n70 );
nand ( n2147, n31, n55 );
xor ( n2148, n25, n36 );
nand ( n2149, n5, n129 );
and ( n2150, n38, n77 );
and ( n2151, n78, n143 );
and ( n2152, n29, n66 );
nor ( n2153, n118, n122 );
and ( n2154, n6, n54 );
nand ( n2155, n11, n56 );
nor ( n2156, n3, n105 );
xor ( n2157, n66, n82 );
nor ( n2158, n61, n136 );
xor ( n2159, n113, n118 );
and ( n2160, n60, n62 );
nor ( n2161, n18, n32 );
xor ( n2162, n4, n28 );
nand ( n2163, n30, n33 );
xor ( n2164, n105, n111 );
nand ( n2165, n102, n113 );
or ( n2166, n52, n141 );
xor ( n2167, n56, n98 );
and ( n2168, n18, n38 );
nand ( n2169, n110, n128 );
or ( n2170, n81, n96 );
and ( n2171, n60, n110 );
nand ( n2172, n40, n63 );
and ( n2173, n33, n74 );
or ( n2174, n34, n106 );
or ( n2175, n85, n137 );
or ( n2176, n27, n57 );
nor ( n2177, n19, n77 );
and ( n2178, n18, n140 );
nor ( n2179, n5, n29 );
nor ( n2180, n21, n130 );
or ( n2181, n13, n121 );
xor ( n2182, n44, n69 );
nor ( n2183, n56, n120 );
xor ( n2184, n34, n55 );
nor ( n2185, n72, n143 );
nand ( n2186, n59, n110 );
nand ( n2187, n44, n98 );
or ( n2188, n64, n140 );
and ( n2189, n79, n111 );
nor ( n2190, n87, n137 );
nand ( n2191, n40, n128 );
xor ( n2192, n44, n52 );
or ( n2193, n31, n103 );
or ( n2194, n33, n55 );
nand ( n2195, n60, n86 );
nand ( n2196, n66, n98 );
xor ( n2197, n57, n139 );
or ( n2198, n3, n70 );
and ( n2199, n12, n131 );
and ( n2200, n29, n53 );
or ( n2201, n73, n88 );
and ( n2202, n21, n28 );
and ( n2203, n7, n65 );
nand ( n2204, n113, n127 );
nor ( n2205, n26, n139 );
xor ( n2206, n92, n117 );
nor ( n2207, n12, n101 );
and ( n2208, n24, n118 );
or ( n2209, n19, n54 );
xor ( n2210, n73, n111 );
nand ( n2211, n29, n126 );
xor ( n2212, n16, n35 );
or ( n2213, n109, n121 );
nor ( n2214, n0, n29 );
and ( n2215, n65, n89 );
xor ( n2216, n64, n142 );
nand ( n2217, n69, n70 );
and ( n2218, n39, n64 );
nor ( n2219, n103, n130 );
xor ( n2220, n107, n126 );
or ( n2221, n120, n134 );
and ( n2222, n41, n120 );
or ( n2223, n69, n97 );
nor ( n2224, n118, n130 );
or ( n2225, n1, n55 );
xor ( n2226, n36, n56 );
xor ( n2227, n20, n130 );
xor ( n2228, n69, n117 );
xor ( n2229, n11, n58 );
nand ( n2230, n35, n87 );
nor ( n2231, n5, n7 );
nor ( n2232, n63, n113 );
nor ( n2233, n22, n69 );
nand ( n2234, n11, n41 );
or ( n2235, n44, n63 );
nand ( n2236, n40, n88 );
nor ( n2237, n42, n111 );
or ( n2238, n30, n80 );
nand ( n2239, n28, n96 );
xor ( n2240, n48, n120 );
xor ( n2241, n94, n129 );
nor ( n2242, n16, n44 );
and ( n2243, n3, n35 );
nand ( n2244, n135, n143 );
nand ( n2245, n91, n137 );
or ( n2246, n11, n134 );
and ( n2247, n11, n130 );
or ( n2248, n25, n112 );
xor ( n2249, n13, n26 );
or ( n2250, n69, n94 );
or ( n2251, n2, n73 );
or ( n2252, n122, n131 );
nand ( n2253, n67, n99 );
nor ( n2254, n86, n87 );
and ( n2255, n27, n87 );
nor ( n2256, n81, n118 );
and ( n2257, n92, n139 );
and ( n2258, n9, n14 );
and ( n2259, n36, n98 );
xor ( n2260, n88, n137 );
xor ( n2261, n116, n132 );
nand ( n2262, n39, n43 );
or ( n2263, n26, n141 );
and ( n2264, n92, n111 );
and ( n2265, n31, n122 );
and ( n2266, n72, n139 );
or ( n2267, n30, n46 );
xor ( n2268, n81, n116 );
nand ( n2269, n18, n22 );
and ( n2270, n83, n133 );
nor ( n2271, n75, n84 );
nand ( n2272, n15, n88 );
or ( n2273, n90, n143 );
or ( n2274, n32, n134 );
or ( n2275, n7, n20 );
or ( n2276, n108, n135 );
and ( n2277, n49, n58 );
xor ( n2278, n103, n104 );
xor ( n2279, n46, n103 );
or ( n2280, n77, n120 );
nor ( n2281, n54, n120 );
xor ( n2282, n14, n88 );
or ( n2283, n70, n140 );
xor ( n2284, n99, n113 );
nor ( n2285, n91, n143 );
and ( n2286, n32, n100 );
nand ( n2287, n91, n123 );
xor ( n2288, n16, n17 );
nor ( n2289, n76, n92 );
or ( n2290, n118, n125 );
and ( n2291, n96, n143 );
nor ( n2292, n88, n98 );
nor ( n2293, n23, n55 );
or ( n2294, n17, n128 );
nor ( n2295, n23, n130 );
or ( n2296, n93, n123 );
nor ( n2297, n0, n3 );
or ( n2298, n4, n113 );
or ( n2299, n7, n51 );
or ( n2300, n8, n45 );
or ( n2301, n68, n70 );
and ( n2302, n66, n95 );
nor ( n2303, n27, n59 );
xor ( n2304, n37, n140 );
and ( n2305, n4, n69 );
nand ( n2306, n59, n126 );
xor ( n2307, n33, n118 );
and ( n2308, n38, n40 );
xor ( n2309, n70, n89 );
xor ( n2310, n68, n104 );
nand ( n2311, n4, n89 );
or ( n2312, n19, n23 );
xor ( n2313, n6, n108 );
nand ( n2314, n68, n125 );
or ( n2315, n57, n79 );
or ( n2316, n38, n115 );
xor ( n2317, n56, n62 );
xor ( n2318, n95, n102 );
or ( n2319, n32, n52 );
nand ( n2320, n73, n125 );
nand ( n2321, n0, n119 );
nor ( n2322, n0, n16 );
nand ( n2323, n66, n114 );
nand ( n2324, n46, n101 );
xor ( n2325, n34, n48 );
nor ( n2326, n92, n121 );
nand ( n2327, n21, n82 );
or ( n2328, n76, n107 );
nand ( n2329, n44, n78 );
and ( n2330, n42, n62 );
or ( n2331, n38, n83 );
and ( n2332, n67, n142 );
nand ( n2333, n24, n49 );
xor ( n2334, n29, n76 );
nand ( n2335, n87, n106 );
xor ( n2336, n26, n137 );
or ( n2337, n43, n91 );
xor ( n2338, n84, n131 );
or ( n2339, n47, n91 );
or ( n2340, n57, n85 );
nor ( n2341, n39, n98 );
nor ( n2342, n4, n105 );
nor ( n2343, n28, n94 );
nor ( n2344, n124, n137 );
xor ( n2345, n64, n69 );
nand ( n2346, n20, n135 );
xor ( n2347, n100, n135 );
xor ( n2348, n93, n113 );
nor ( n2349, n3, n50 );
and ( n2350, n118, n123 );
nor ( n2351, n79, n82 );
or ( n2352, n78, n105 );
nand ( n2353, n12, n24 );
and ( n2354, n10, n71 );
nand ( n2355, n112, n143 );
or ( n2356, n21, n120 );
xor ( n2357, n34, n67 );
and ( n2358, n81, n91 );
xor ( n2359, n86, n134 );
nor ( n2360, n23, n34 );
nor ( n2361, n133, n142 );
and ( n2362, n13, n25 );
nand ( n2363, n87, n120 );
xor ( n2364, n68, n69 );
xor ( n2365, n101, n103 );
nand ( n2366, n10, n78 );
or ( n2367, n66, n68 );
or ( n2368, n0, n108 );
and ( n2369, n105, n109 );
or ( n2370, n55, n56 );
nand ( n2371, n17, n96 );
and ( n2372, n52, n120 );
or ( n2373, n71, n101 );
or ( n2374, n10, n15 );
nand ( n2375, n4, n117 );
nor ( n2376, n86, n97 );
nand ( n2377, n10, n115 );
nand ( n2378, n11, n79 );
or ( n2379, n56, n104 );
nand ( n2380, n34, n117 );
xor ( n2381, n19, n121 );
or ( n2382, n29, n108 );
and ( n2383, n115, n142 );
and ( n2384, n59, n94 );
nand ( n2385, n15, n91 );
xor ( n2386, n15, n43 );
or ( n2387, n62, n73 );
and ( n2388, n89, n96 );
and ( n2389, n49, n94 );
nand ( n2390, n95, n110 );
xor ( n2391, n16, n38 );
or ( n2392, n22, n64 );
nand ( n2393, n27, n103 );
xor ( n2394, n10, n49 );
nor ( n2395, n10, n28 );
nand ( n2396, n76, n115 );
nand ( n2397, n19, n84 );
nand ( n2398, n90, n104 );
xor ( n2399, n36, n138 );
nand ( n2400, n18, n24 );
or ( n2401, n2, n114 );
nor ( n2402, n71, n135 );
or ( n2403, n67, n87 );
nand ( n2404, n52, n74 );
and ( n2405, n52, n102 );
and ( n2406, n48, n50 );
or ( n2407, n22, n32 );
and ( n2408, n77, n88 );
xor ( n2409, n69, n126 );
or ( n2410, n8, n23 );
and ( n2411, n63, n73 );
or ( n2412, n93, n94 );
nand ( n2413, n29, n70 );
or ( n2414, n63, n64 );
xor ( n2415, n60, n141 );
nor ( n2416, n24, n101 );
and ( n2417, n94, n109 );
nor ( n2418, n2, n56 );
nor ( n2419, n1, n14 );
nand ( n2420, n3, n69 );
xor ( n2421, n10, n34 );
nand ( n2422, n53, n128 );
xor ( n2423, n48, n56 );
and ( n2424, n113, n140 );
and ( n2425, n21, n122 );
xor ( n2426, n55, n80 );
or ( n2427, n4, n27 );
xor ( n2428, n51, n113 );
xor ( n2429, n9, n33 );
xor ( n2430, n33, n99 );
and ( n2431, n28, n120 );
or ( n2432, n26, n45 );
nor ( n2433, n44, n139 );
nor ( n2434, n96, n121 );
nor ( n2435, n58, n74 );
or ( n2436, n112, n129 );
nor ( n2437, n3, n103 );
xor ( n2438, n92, n131 );
nand ( n2439, n72, n89 );
nor ( n2440, n22, n85 );
and ( n2441, n6, n77 );
or ( n2442, n62, n77 );
nor ( n2443, n10, n23 );
or ( n2444, n0, n7 );
nand ( n2445, n48, n80 );
or ( n2446, n45, n46 );
or ( n2447, n73, n113 );
and ( n2448, n49, n130 );
nand ( n2449, n112, n125 );
nand ( n2450, n18, n109 );
or ( n2451, n128, n143 );
and ( n2452, n54, n121 );
xor ( n2453, n60, n124 );
nand ( n2454, n1, n135 );
and ( n2455, n71, n102 );
or ( n2456, n5, n113 );
and ( n2457, n95, n119 );
or ( n2458, n34, n143 );
nand ( n2459, n58, n67 );
xor ( n2460, n111, n112 );
nand ( n2461, n23, n88 );
nand ( n2462, n47, n67 );
or ( n2463, n33, n106 );
nor ( n2464, n29, n50 );
nor ( n2465, n26, n65 );
or ( n2466, n48, n86 );
or ( n2467, n26, n110 );
nor ( n2468, n51, n107 );
nand ( n2469, n9, n80 );
or ( n2470, n16, n102 );
and ( n2471, n1, n65 );
nand ( n2472, n42, n135 );
nor ( n2473, n24, n81 );
and ( n2474, n54, n93 );
nand ( n2475, n6, n26 );
and ( n2476, n36, n84 );
nand ( n2477, n115, n140 );
or ( n2478, n102, n112 );
or ( n2479, n104, n141 );
and ( n2480, n7, n34 );
or ( n2481, n11, n91 );
nor ( n2482, n49, n72 );
xor ( n2483, n60, n82 );
nand ( n2484, n91, n109 );
or ( n2485, n46, n54 );
nor ( n2486, n62, n78 );
xor ( n2487, n11, n126 );
nand ( n2488, n20, n30 );
nor ( n2489, n43, n45 );
and ( n2490, n17, n111 );
xor ( n2491, n54, n79 );
nor ( n2492, n87, n112 );
nand ( n2493, n121, n136 );
xor ( n2494, n121, n142 );
xor ( n2495, n87, n101 );
and ( n2496, n31, n34 );
and ( n2497, n10, n111 );
or ( n2498, n112, n139 );
or ( n2499, n137, n139 );
xor ( n2500, n45, n121 );
nand ( n2501, n34, n130 );
and ( n2502, n38, n86 );
nand ( n2503, n19, n105 );
xor ( n2504, n10, n65 );
xor ( n2505, n88, n104 );
and ( n2506, n2, n19 );
nand ( n2507, n0, n78 );
nor ( n2508, n34, n72 );
nor ( n2509, n6, n45 );
xor ( n2510, n38, n94 );
and ( n2511, n35, n135 );
nor ( n2512, n8, n57 );
xor ( n2513, n41, n112 );
nor ( n2514, n21, n26 );
and ( n2515, n3, n31 );
nor ( n2516, n77, n101 );
nand ( n2517, n111, n130 );
nor ( n2518, n14, n70 );
or ( n2519, n41, n63 );
nor ( n2520, n60, n132 );
xor ( n2521, n23, n113 );
nand ( n2522, n17, n88 );
nor ( n2523, n22, n33 );
nor ( n2524, n53, n134 );
nor ( n2525, n127, n139 );
nor ( n2526, n13, n91 );
nand ( n2527, n22, n112 );
nand ( n2528, n54, n74 );
and ( n2529, n48, n55 );
nand ( n2530, n83, n84 );
nand ( n2531, n14, n84 );
or ( n2532, n36, n87 );
or ( n2533, n62, n122 );
nand ( n2534, n34, n109 );
xor ( n2535, n79, n106 );
xor ( n2536, n19, n55 );
and ( n2537, n19, n123 );
nand ( n2538, n68, n76 );
nand ( n2539, n74, n86 );
xor ( n2540, n92, n140 );
xor ( n2541, n11, n31 );
nand ( n2542, n3, n72 );
xor ( n2543, n96, n126 );
xor ( n2544, n35, n127 );
nand ( n2545, n67, n85 );
or ( n2546, n42, n118 );
nor ( n2547, n40, n129 );
xor ( n2548, n78, n80 );
or ( n2549, n34, n134 );
xor ( n2550, n17, n77 );
nor ( n2551, n56, n136 );
or ( n2552, n54, n101 );
nand ( n2553, n30, n126 );
nand ( n2554, n62, n101 );
xor ( n2555, n3, n65 );
xor ( n2556, n22, n122 );
nand ( n2557, n15, n118 );
nand ( n2558, n62, n107 );
nand ( n2559, n1, n22 );
and ( n2560, n94, n114 );
and ( n2561, n20, n72 );
nor ( n2562, n19, n135 );
or ( n2563, n51, n84 );
nand ( n2564, n80, n116 );
or ( n2565, n4, n124 );
xor ( n2566, n1, n107 );
nand ( n2567, n3, n82 );
nand ( n2568, n46, n92 );
and ( n2569, n31, n41 );
xor ( n2570, n74, n102 );
nor ( n2571, n130, n140 );
nand ( n2572, n48, n99 );
xor ( n2573, n85, n118 );
xor ( n2574, n64, n136 );
xor ( n2575, n48, n58 );
nand ( n2576, n42, n55 );
and ( n2577, n102, n141 );
nand ( n2578, n23, n124 );
nor ( n2579, n21, n129 );
nand ( n2580, n75, n113 );
nand ( n2581, n18, n129 );
xor ( n2582, n77, n80 );
or ( n2583, n122, n142 );
nand ( n2584, n44, n80 );
or ( n2585, n19, n101 );
or ( n2586, n8, n90 );
nand ( n2587, n41, n119 );
and ( n2588, n65, n121 );
nor ( n2589, n15, n102 );
nand ( n2590, n99, n126 );
xor ( n2591, n65, n112 );
nor ( n2592, n7, n100 );
and ( n2593, n14, n54 );
nand ( n2594, n66, n127 );
xor ( n2595, n52, n75 );
xor ( n2596, n0, n99 );
nand ( n2597, n117, n119 );
or ( n2598, n6, n57 );
nor ( n2599, n12, n137 );
or ( n2600, n9, n24 );
nor ( n2601, n4, n140 );
xor ( n2602, n46, n56 );
nor ( n2603, n42, n107 );
nand ( n2604, n106, n109 );
nand ( n2605, n8, n9 );
xor ( n2606, n70, n84 );
xor ( n2607, n49, n140 );
nand ( n2608, n83, n138 );
and ( n2609, n80, n94 );
and ( n2610, n28, n89 );
xor ( n2611, n33, n94 );
xor ( n2612, n64, n101 );
and ( n2613, n52, n62 );
or ( n2614, n42, n127 );
xor ( n2615, n8, n15 );
nor ( n2616, n56, n59 );
or ( n2617, n131, n139 );
nand ( n2618, n116, n143 );
and ( n2619, n57, n135 );
nor ( n2620, n13, n51 );
or ( n2621, n43, n89 );
or ( n2622, n57, n69 );
nand ( n2623, n99, n121 );
xor ( n2624, n15, n85 );
nand ( n2625, n101, n127 );
xor ( n2626, n76, n119 );
nand ( n2627, n53, n111 );
and ( n2628, n75, n127 );
xor ( n2629, n57, n95 );
and ( n2630, n23, n138 );
nor ( n2631, n43, n114 );
nand ( n2632, n3, n60 );
or ( n2633, n28, n62 );
nor ( n2634, n48, n135 );
nand ( n2635, n18, n83 );
nor ( n2636, n19, n89 );
xor ( n2637, n9, n43 );
nor ( n2638, n39, n59 );
and ( n2639, n57, n90 );
nor ( n2640, n52, n60 );
xor ( n2641, n14, n104 );
xor ( n2642, n35, n143 );
and ( n2643, n130, n135 );
or ( n2644, n32, n121 );
and ( n2645, n77, n115 );
and ( n2646, n136, n139 );
or ( n2647, n83, n118 );
and ( n2648, n52, n132 );
nor ( n2649, n23, n73 );
nor ( n2650, n9, n108 );
nand ( n2651, n45, n125 );
and ( n2652, n23, n85 );
xor ( n2653, n120, n126 );
nand ( n2654, n26, n34 );
or ( n2655, n99, n112 );
or ( n2656, n9, n142 );
nor ( n2657, n85, n102 );
or ( n2658, n5, n65 );
nand ( n2659, n2, n121 );
and ( n2660, n8, n109 );
xor ( n2661, n63, n76 );
and ( n2662, n3, n132 );
or ( n2663, n36, n69 );
and ( n2664, n25, n93 );
and ( n2665, n79, n132 );
nor ( n2666, n42, n99 );
or ( n2667, n60, n72 );
nand ( n2668, n137, n142 );
and ( n2669, n107, n120 );
xor ( n2670, n51, n88 );
nor ( n2671, n117, n127 );
xor ( n2672, n12, n43 );
nand ( n2673, n12, n15 );
or ( n2674, n96, n106 );
xor ( n2675, n22, n79 );
nor ( n2676, n64, n119 );
nor ( n2677, n23, n82 );
nand ( n2678, n18, n54 );
nor ( n2679, n124, n129 );
and ( n2680, n70, n114 );
nand ( n2681, n4, n136 );
nor ( n2682, n30, n114 );
and ( n2683, n35, n141 );
nand ( n2684, n70, n112 );
or ( n2685, n19, n98 );
or ( n2686, n5, n44 );
or ( n2687, n51, n65 );
or ( n2688, n89, n143 );
xor ( n2689, n5, n120 );
or ( n2690, n80, n136 );
and ( n2691, n8, n76 );
or ( n2692, n36, n94 );
and ( n2693, n23, n96 );
xor ( n2694, n81, n105 );
or ( n2695, n8, n58 );
nor ( n2696, n43, n112 );
and ( n2697, n71, n108 );
nor ( n2698, n66, n96 );
nand ( n2699, n110, n133 );
nor ( n2700, n62, n94 );
xor ( n2701, n13, n135 );
nor ( n2702, n53, n124 );
and ( n2703, n18, n139 );
and ( n2704, n55, n58 );
nand ( n2705, n124, n134 );
and ( n2706, n44, n77 );
and ( n2707, n11, n22 );
nand ( n2708, n60, n77 );
and ( n2709, n14, n76 );
nand ( n2710, n53, n79 );
or ( n2711, n0, n82 );
nand ( n2712, n83, n113 );
nor ( n2713, n23, n108 );
xor ( n2714, n19, n78 );
nand ( n2715, n16, n93 );
nor ( n2716, n9, n110 );
nand ( n2717, n61, n95 );
nor ( n2718, n9, n76 );
and ( n2719, n107, n115 );
nand ( n2720, n92, n129 );
xor ( n2721, n42, n59 );
and ( n2722, n93, n135 );
xor ( n2723, n8, n87 );
nand ( n2724, n99, n115 );
nand ( n2725, n35, n103 );
and ( n2726, n4, n82 );
and ( n2727, n49, n117 );
and ( n2728, n29, n132 );
and ( n2729, n24, n79 );
nand ( n2730, n34, n98 );
and ( n2731, n90, n121 );
xor ( n2732, n18, n123 );
and ( n2733, n44, n49 );
or ( n2734, n38, n51 );
or ( n2735, n31, n113 );
or ( n2736, n64, n109 );
xor ( n2737, n41, n74 );
or ( n2738, n48, n103 );
and ( n2739, n119, n140 );
nor ( n2740, n48, n104 );
or ( n2741, n22, n123 );
and ( n2742, n38, n129 );
nand ( n2743, n63, n72 );
or ( n2744, n89, n118 );
nand ( n2745, n27, n35 );
xor ( n2746, n53, n106 );
nor ( n2747, n26, n42 );
and ( n2748, n112, n132 );
or ( n2749, n40, n48 );
and ( n2750, n55, n126 );
nor ( n2751, n37, n133 );
nor ( n2752, n59, n72 );
xor ( n2753, n37, n107 );
and ( n2754, n77, n122 );
nand ( n2755, n36, n123 );
and ( n2756, n29, n47 );
nand ( n2757, n51, n129 );
xor ( n2758, n12, n103 );
nor ( n2759, n105, n138 );
and ( n2760, n30, n96 );
nand ( n2761, n21, n45 );
xor ( n2762, n107, n111 );
nand ( n2763, n49, n111 );
nor ( n2764, n69, n106 );
nor ( n2765, n85, n127 );
or ( n2766, n37, n81 );
nor ( n2767, n128, n137 );
nand ( n2768, n80, n106 );
xor ( n2769, n71, n99 );
and ( n2770, n117, n124 );
nor ( n2771, n24, n87 );
xor ( n2772, n51, n100 );
or ( n2773, n10, n90 );
xor ( n2774, n30, n81 );
and ( n2775, n0, n23 );
and ( n2776, n36, n77 );
nor ( n2777, n38, n63 );
and ( n2778, n14, n71 );
nor ( n2779, n89, n105 );
or ( n2780, n59, n80 );
nor ( n2781, n90, n134 );
and ( n2782, n20, n76 );
or ( n2783, n16, n135 );
xor ( n2784, n92, n103 );
xor ( n2785, n20, n29 );
xor ( n2786, n22, n55 );
nor ( n2787, n54, n99 );
nor ( n2788, n21, n47 );
or ( n2789, n66, n115 );
xor ( n2790, n92, n105 );
nand ( n2791, n43, n76 );
nand ( n2792, n24, n96 );
or ( n2793, n82, n106 );
nor ( n2794, n38, n48 );
or ( n2795, n32, n85 );
and ( n2796, n16, n134 );
or ( n2797, n24, n141 );
and ( n2798, n68, n90 );
or ( n2799, n90, n141 );
xor ( n2800, n80, n101 );
nand ( n2801, n50, n129 );
nor ( n2802, n6, n119 );
or ( n2803, n53, n58 );
and ( n2804, n98, n120 );
nor ( n2805, n130, n139 );
or ( n2806, n12, n70 );
xor ( n2807, n0, n134 );
nor ( n2808, n87, n111 );
nor ( n2809, n50, n81 );
nor ( n2810, n69, n132 );
nand ( n2811, n83, n96 );
and ( n2812, n10, n47 );
nand ( n2813, n71, n132 );
xor ( n2814, n0, n109 );
and ( n2815, n53, n90 );
xor ( n2816, n31, n72 );
and ( n2817, n107, n139 );
nor ( n2818, n26, n73 );
nor ( n2819, n20, n134 );
nand ( n2820, n58, n125 );
nand ( n2821, n35, n38 );
and ( n2822, n95, n122 );
nand ( n2823, n23, n142 );
or ( n2824, n49, n57 );
and ( n2825, n129, n140 );
and ( n2826, n1, n58 );
xor ( n2827, n92, n112 );
nand ( n2828, n61, n115 );
nand ( n2829, n0, n67 );
xor ( n2830, n36, n71 );
and ( n2831, n20, n107 );
or ( n2832, n32, n135 );
and ( n2833, n12, n90 );
xor ( n2834, n27, n130 );
and ( n2835, n18, n46 );
and ( n2836, n92, n109 );
or ( n2837, n20, n21 );
and ( n2838, n35, n104 );
xor ( n2839, n10, n127 );
xor ( n2840, n13, n133 );
and ( n2841, n17, n37 );
nor ( n2842, n97, n140 );
nand ( n2843, n35, n130 );
and ( n2844, n22, n81 );
nor ( n2845, n89, n141 );
and ( n2846, n96, n133 );
and ( n2847, n22, n116 );
or ( n2848, n5, n79 );
xor ( n2849, n80, n142 );
nand ( n2850, n76, n85 );
nand ( n2851, n33, n125 );
xor ( n2852, n80, n134 );
nor ( n2853, n11, n72 );
and ( n2854, n111, n119 );
or ( n2855, n6, n94 );
nand ( n2856, n66, n110 );
xor ( n2857, n20, n47 );
nor ( n2858, n82, n99 );
xor ( n2859, n4, n61 );
xor ( n2860, n55, n63 );
nor ( n2861, n8, n125 );
xor ( n2862, n9, n40 );
or ( n2863, n41, n66 );
and ( n2864, n87, n118 );
and ( n2865, n103, n127 );
and ( n2866, n4, n35 );
or ( n2867, n87, n129 );
xor ( n2868, n40, n108 );
xor ( n2869, n118, n142 );
xor ( n2870, n24, n43 );
and ( n2871, n5, n95 );
nor ( n2872, n38, n97 );
nor ( n2873, n63, n82 );
nand ( n2874, n18, n56 );
xor ( n2875, n3, n48 );
nor ( n2876, n15, n99 );
xor ( n2877, n113, n137 );
xor ( n2878, n19, n126 );
nand ( n2879, n8, n56 );
nor ( n2880, n45, n86 );
or ( n2881, n51, n71 );
or ( n2882, n21, n105 );
xor ( n2883, n53, n138 );
or ( n2884, n71, n85 );
nand ( n2885, n27, n93 );
nand ( n2886, n16, n20 );
xor ( n2887, n67, n140 );
xor ( n2888, n8, n128 );
xor ( n2889, n12, n138 );
nor ( n2890, n56, n119 );
nand ( n2891, n46, n102 );
nor ( n2892, n111, n124 );
or ( n2893, n24, n54 );
nor ( n2894, n42, n45 );
or ( n2895, n21, n117 );
nand ( n2896, n6, n103 );
nor ( n2897, n38, n44 );
and ( n2898, n73, n84 );
xor ( n2899, n21, n66 );
xor ( n2900, n78, n130 );
nand ( n2901, n45, n104 );
nand ( n2902, n62, n121 );
and ( n2903, n62, n134 );
or ( n2904, n29, n112 );
and ( n2905, n80, n85 );
nor ( n2906, n11, n75 );
nand ( n2907, n7, n129 );
and ( n2908, n4, n123 );
or ( n2909, n82, n130 );
and ( n2910, n18, n57 );
xor ( n2911, n40, n60 );
or ( n2912, n22, n76 );
and ( n2913, n63, n99 );
and ( n2914, n108, n111 );
and ( n2915, n75, n136 );
nand ( n2916, n45, n120 );
or ( n2917, n27, n61 );
or ( n2918, n109, n131 );
or ( n2919, n4, n65 );
nand ( n2920, n10, n22 );
or ( n2921, n1, n106 );
and ( n2922, n100, n133 );
and ( n2923, n33, n136 );
nor ( n2924, n63, n136 );
or ( n2925, n58, n94 );
and ( n2926, n76, n99 );
or ( n2927, n38, n92 );
and ( n2928, n7, n74 );
or ( n2929, n8, n53 );
nand ( n2930, n18, n131 );
and ( n2931, n93, n139 );
nor ( n2932, n90, n128 );
xor ( n2933, n13, n63 );
nor ( n2934, n4, n56 );
nand ( n2935, n29, n139 );
or ( n2936, n15, n73 );
nor ( n2937, n17, n136 );
and ( n2938, n104, n130 );
nor ( n2939, n30, n73 );
and ( n2940, n25, n103 );
xor ( n2941, n27, n37 );
or ( n2942, n28, n123 );
nor ( n2943, n85, n134 );
nand ( n2944, n51, n90 );
and ( n2945, n105, n133 );
nand ( n2946, n15, n83 );
or ( n2947, n48, n108 );
xor ( n2948, n52, n83 );
or ( n2949, n26, n74 );
xor ( n2950, n10, n69 );
xor ( n2951, n64, n89 );
nand ( n2952, n46, n84 );
nand ( n2953, n30, n42 );
nand ( n2954, n54, n113 );
and ( n2955, n66, n123 );
nand ( n2956, n73, n140 );
or ( n2957, n26, n140 );
or ( n2958, n2, n96 );
and ( n2959, n77, n89 );
nor ( n2960, n92, n98 );
xor ( n2961, n85, n123 );
and ( n2962, n69, n100 );
nor ( n2963, n15, n22 );
and ( n2964, n44, n83 );
or ( n2965, n58, n102 );
and ( n2966, n37, n109 );
or ( n2967, n6, n136 );
nor ( n2968, n2, n31 );
and ( n2969, n9, n51 );
and ( n2970, n125, n137 );
xor ( n2971, n32, n122 );
and ( n2972, n85, n124 );
nor ( n2973, n81, n100 );
nor ( n2974, n46, n134 );
and ( n2975, n111, n133 );
nor ( n2976, n14, n44 );
and ( n2977, n61, n63 );
nand ( n2978, n29, n120 );
nand ( n2979, n68, n84 );
and ( n2980, n121, n125 );
nor ( n2981, n59, n106 );
nand ( n2982, n7, n32 );
nor ( n2983, n93, n120 );
nor ( n2984, n38, n112 );
or ( n2985, n112, n114 );
or ( n2986, n87, n121 );
and ( n2987, n21, n100 );
nand ( n2988, n56, n100 );
or ( n2989, n96, n102 );
nand ( n2990, n55, n74 );
xor ( n2991, n34, n82 );
nor ( n2992, n81, n89 );
or ( n2993, n123, n135 );
or ( n2994, n14, n134 );
or ( n2995, n88, n107 );
nand ( n2996, n34, n113 );
and ( n2997, n32, n86 );
nor ( n2998, n8, n71 );
nor ( n2999, n99, n142 );
nand ( n3000, n29, n113 );
or ( n3001, n5, n78 );
or ( n3002, n115, n133 );
nand ( n3003, n5, n106 );
or ( n3004, n111, n113 );
nor ( n3005, n64, n139 );
or ( n3006, n108, n126 );
nor ( n3007, n29, n86 );
nor ( n3008, n13, n31 );
or ( n3009, n71, n138 );
or ( n3010, n20, n131 );
nand ( n3011, n85, n110 );
or ( n3012, n1, n32 );
or ( n3013, n92, n110 );
xor ( n3014, n38, n105 );
and ( n3015, n14, n79 );
or ( n3016, n2, n40 );
xor ( n3017, n93, n99 );
xor ( n3018, n38, n126 );
nor ( n3019, n72, n82 );
nand ( n3020, n46, n57 );
or ( n3021, n8, n96 );
nand ( n3022, n40, n141 );
or ( n3023, n78, n103 );
nand ( n3024, n35, n55 );
nor ( n3025, n8, n25 );
xor ( n3026, n2, n90 );
xor ( n3027, n31, n46 );
and ( n3028, n73, n110 );
and ( n3029, n56, n82 );
xor ( n3030, n98, n124 );
xor ( n3031, n36, n126 );
and ( n3032, n68, n122 );
and ( n3033, n45, n70 );
nor ( n3034, n23, n98 );
or ( n3035, n53, n103 );
and ( n3036, n7, n33 );
nand ( n3037, n2, n116 );
nor ( n3038, n10, n45 );
nand ( n3039, n7, n69 );
or ( n3040, n58, n121 );
and ( n3041, n119, n143 );
xor ( n3042, n69, n108 );
xor ( n3043, n10, n38 );
and ( n3044, n89, n124 );
nor ( n3045, n61, n78 );
xor ( n3046, n77, n104 );
nand ( n3047, n126, n143 );
and ( n3048, n37, n47 );
xor ( n3049, n106, n116 );
nor ( n3050, n27, n85 );
nand ( n3051, n24, n77 );
nand ( n3052, n30, n110 );
nand ( n3053, n47, n98 );
nand ( n3054, n80, n132 );
and ( n3055, n3, n49 );
or ( n3056, n23, n128 );
nor ( n3057, n53, n130 );
nor ( n3058, n14, n27 );
and ( n3059, n22, n30 );
or ( n3060, n10, n27 );
and ( n3061, n14, n80 );
xor ( n3062, n17, n79 );
nand ( n3063, n1, n8 );
xor ( n3064, n96, n104 );
nand ( n3065, n9, n126 );
and ( n3066, n41, n44 );
nor ( n3067, n75, n92 );
nor ( n3068, n24, n135 );
or ( n3069, n4, n91 );
nand ( n3070, n37, n116 );
or ( n3071, n103, n108 );
nor ( n3072, n109, n124 );
and ( n3073, n42, n66 );
and ( n3074, n85, n98 );
xor ( n3075, n32, n93 );
and ( n3076, n32, n88 );
and ( n3077, n61, n80 );
nand ( n3078, n96, n142 );
or ( n3079, n55, n102 );
or ( n3080, n34, n104 );
and ( n3081, n3, n73 );
and ( n3082, n49, n68 );
or ( n3083, n31, n42 );
and ( n3084, n45, n137 );
or ( n3085, n114, n135 );
nor ( n3086, n25, n62 );
and ( n3087, n6, n116 );
or ( n3088, n57, n114 );
or ( n3089, n79, n113 );
or ( n3090, n67, n111 );
nand ( n3091, n100, n125 );
nor ( n3092, n37, n96 );
nor ( n3093, n49, n107 );
and ( n3094, n26, n27 );
or ( n3095, n36, n110 );
and ( n3096, n117, n118 );
and ( n3097, n31, n110 );
or ( n3098, n36, n68 );
and ( n3099, n86, n135 );
xor ( n3100, n11, n139 );
or ( n3101, n73, n119 );
xor ( n3102, n113, n119 );
or ( n3103, n11, n135 );
or ( n3104, n44, n45 );
or ( n3105, n11, n37 );
and ( n3106, n65, n115 );
and ( n3107, n104, n113 );
and ( n3108, n3, n98 );
or ( n3109, n27, n67 );
nor ( n3110, n10, n125 );
or ( n3111, n60, n78 );
nor ( n3112, n30, n64 );
xor ( n3113, n37, n126 );
nand ( n3114, n14, n128 );
nand ( n3115, n32, n68 );
and ( n3116, n0, n22 );
xor ( n3117, n12, n18 );
nand ( n3118, n114, n121 );
nor ( n3119, n21, n75 );
and ( n3120, n104, n124 );
xor ( n3121, n135, n136 );
xor ( n3122, n50, n53 );
xor ( n3123, n61, n97 );
or ( n3124, n19, n74 );
nand ( n3125, n17, n47 );
and ( n3126, n17, n33 );
or ( n3127, n33, n133 );
nand ( n3128, n11, n90 );
nand ( n3129, n18, n77 );
nand ( n3130, n16, n74 );
and ( n3131, n72, n105 );
nand ( n3132, n72, n84 );
nand ( n3133, n15, n139 );
nand ( n3134, n11, n53 );
or ( n3135, n10, n41 );
and ( n3136, n16, n41 );
nor ( n3137, n98, n142 );
xor ( n3138, n89, n125 );
and ( n3139, n71, n103 );
xor ( n3140, n19, n79 );
nor ( n3141, n67, n77 );
xor ( n3142, n30, n92 );
or ( n3143, n6, n18 );
nor ( n3144, n15, n92 );
and ( n3145, n88, n120 );
nor ( n3146, n118, n124 );
nor ( n3147, n35, n122 );
or ( n3148, n46, n79 );
or ( n3149, n21, n41 );
nand ( n3150, n7, n42 );
nor ( n3151, n22, n101 );
nand ( n3152, n95, n139 );
nand ( n3153, n69, n116 );
nor ( n3154, n31, n117 );
nand ( n3155, n65, n127 );
nand ( n3156, n115, n121 );
nor ( n3157, n84, n119 );
nand ( n3158, n26, n72 );
nand ( n3159, n126, n131 );
or ( n3160, n16, n58 );
nor ( n3161, n8, n138 );
nand ( n3162, n64, n143 );
nor ( n3163, n7, n84 );
xor ( n3164, n23, n60 );
nor ( n3165, n1, n92 );
nor ( n3166, n16, n91 );
nand ( n3167, n60, n76 );
nand ( n3168, n30, n143 );
and ( n3169, n87, n131 );
nor ( n3170, n25, n98 );
or ( n3171, n55, n70 );
or ( n3172, n86, n142 );
and ( n3173, n28, n117 );
nor ( n3174, n6, n127 );
or ( n3175, n57, n137 );
nand ( n3176, n52, n118 );
and ( n3177, n46, n71 );
nor ( n3178, n39, n80 );
nor ( n3179, n84, n132 );
nor ( n3180, n80, n113 );
nor ( n3181, n2, n134 );
xor ( n3182, n5, n43 );
nor ( n3183, n6, n105 );
and ( n3184, n21, n67 );
xor ( n3185, n22, n119 );
xor ( n3186, n7, n54 );
nor ( n3187, n29, n128 );
xor ( n3188, n98, n122 );
nand ( n3189, n2, n112 );
nor ( n3190, n8, n31 );
xor ( n3191, n67, n92 );
xor ( n3192, n108, n132 );
xor ( n3193, n16, n106 );
nor ( n3194, n72, n92 );
nand ( n3195, n96, n138 );
xor ( n3196, n76, n113 );
xor ( n3197, n107, n125 );
nand ( n3198, n1, n71 );
nor ( n3199, n14, n105 );
and ( n3200, n35, n72 );
xor ( n3201, n23, n56 );
nand ( n3202, n40, n139 );
xor ( n3203, n7, n37 );
xor ( n3204, n6, n137 );
nor ( n3205, n7, n47 );
or ( n3206, n26, n129 );
nor ( n3207, n19, n20 );
or ( n3208, n83, n86 );
and ( n3209, n50, n75 );
xor ( n3210, n1, n89 );
xor ( n3211, n75, n119 );
or ( n3212, n49, n136 );
or ( n3213, n71, n133 );
xor ( n3214, n82, n97 );
nand ( n3215, n36, n88 );
nand ( n3216, n34, n139 );
and ( n3217, n80, n105 );
xor ( n3218, n17, n31 );
xor ( n3219, n36, n42 );
nor ( n3220, n44, n138 );
and ( n3221, n0, n79 );
nand ( n3222, n26, n30 );
and ( n3223, n13, n99 );
and ( n3224, n30, n63 );
nand ( n3225, n97, n122 );
or ( n3226, n52, n121 );
nand ( n3227, n35, n94 );
nor ( n3228, n21, n80 );
nor ( n3229, n123, n134 );
nand ( n3230, n89, n128 );
or ( n3231, n18, n63 );
nand ( n3232, n21, n124 );
or ( n3233, n8, n52 );
or ( n3234, n70, n88 );
xor ( n3235, n95, n135 );
xor ( n3236, n31, n63 );
nor ( n3237, n71, n91 );
xor ( n3238, n8, n130 );
and ( n3239, n23, n140 );
or ( n3240, n35, n40 );
or ( n3241, n50, n85 );
nor ( n3242, n53, n73 );
nor ( n3243, n75, n89 );
nor ( n3244, n39, n133 );
and ( n3245, n55, n75 );
or ( n3246, n96, n139 );
nor ( n3247, n103, n106 );
xor ( n3248, n60, n128 );
nand ( n3249, n48, n98 );
or ( n3250, n110, n120 );
xor ( n3251, n22, n65 );
nand ( n3252, n49, n74 );
xor ( n3253, n121, n133 );
nor ( n3254, n16, n118 );
nor ( n3255, n26, n105 );
or ( n3256, n44, n141 );
and ( n3257, n16, n104 );
and ( n3258, n30, n85 );
nor ( n3259, n38, n82 );
or ( n3260, n36, n101 );
or ( n3261, n12, n48 );
xor ( n3262, n94, n125 );
xor ( n3263, n52, n124 );
or ( n3264, n25, n132 );
nand ( n3265, n125, n140 );
nand ( n3266, n35, n96 );
and ( n3267, n98, n107 );
xor ( n3268, n28, n90 );
nor ( n3269, n41, n111 );
xor ( n3270, n64, n94 );
xor ( n3271, n19, n129 );
nand ( n3272, n23, n68 );
nand ( n3273, n114, n134 );
nand ( n3274, n12, n107 );
nand ( n3275, n102, n127 );
xor ( n3276, n7, n63 );
nor ( n3277, n88, n97 );
and ( n3278, n84, n91 );
nor ( n3279, n64, n131 );
nand ( n3280, n73, n83 );
xor ( n3281, n10, n124 );
nor ( n3282, n37, n91 );
xor ( n3283, n23, n100 );
nor ( n3284, n14, n140 );
and ( n3285, n96, n97 );
nand ( n3286, n0, n87 );
or ( n3287, n27, n41 );
xor ( n3288, n9, n132 );
nand ( n3289, n68, n132 );
nand ( n3290, n32, n77 );
xor ( n3291, n70, n115 );
or ( n3292, n13, n81 );
or ( n3293, n34, n97 );
and ( n3294, n38, n104 );
nor ( n3295, n25, n56 );
and ( n3296, n85, n111 );
or ( n3297, n28, n38 );
nand ( n3298, n27, n102 );
or ( n3299, n4, n73 );
or ( n3300, n23, n97 );
or ( n3301, n69, n91 );
nand ( n3302, n56, n110 );
nand ( n3303, n4, n53 );
xor ( n3304, n42, n85 );
and ( n3305, n7, n83 );
nand ( n3306, n85, n99 );
xor ( n3307, n21, n40 );
nor ( n3308, n0, n74 );
nor ( n3309, n54, n55 );
nor ( n3310, n114, n126 );
xor ( n3311, n53, n75 );
and ( n3312, n42, n90 );
or ( n3313, n62, n72 );
nand ( n3314, n14, n142 );
nor ( n3315, n70, n116 );
nand ( n3316, n39, n67 );
and ( n3317, n4, n128 );
nor ( n3318, n86, n104 );
and ( n3319, n54, n89 );
nand ( n3320, n17, n104 );
or ( n3321, n86, n108 );
or ( n3322, n8, n127 );
or ( n3323, n2, n135 );
xor ( n3324, n10, n110 );
xor ( n3325, n8, n88 );
and ( n3326, n132, n134 );
and ( n3327, n41, n50 );
and ( n3328, n5, n62 );
and ( n3329, n24, n89 );
or ( n3330, n126, n139 );
nor ( n3331, n77, n85 );
or ( n3332, n23, n36 );
and ( n3333, n80, n138 );
or ( n3334, n63, n140 );
or ( n3335, n2, n97 );
nor ( n3336, n15, n71 );
nor ( n3337, n101, n132 );
and ( n3338, n93, n108 );
nand ( n3339, n14, n17 );
nand ( n3340, n25, n49 );
and ( n3341, n32, n110 );
nand ( n3342, n37, n61 );
or ( n3343, n40, n99 );
nor ( n3344, n84, n110 );
and ( n3345, n17, n86 );
nor ( n3346, n6, n88 );
and ( n3347, n115, n134 );
and ( n3348, n0, n81 );
or ( n3349, n51, n138 );
nor ( n3350, n94, n140 );
nor ( n3351, n0, n107 );
or ( n3352, n3, n77 );
xor ( n3353, n69, n72 );
nor ( n3354, n43, n116 );
or ( n3355, n35, n93 );
nor ( n3356, n35, n85 );
xor ( n3357, n34, n136 );
xor ( n3358, n69, n86 );
xor ( n3359, n3, n86 );
xor ( n3360, n18, n41 );
nor ( n3361, n59, n60 );
nor ( n3362, n41, n55 );
or ( n3363, n12, n59 );
nand ( n3364, n108, n136 );
xor ( n3365, n125, n133 );
nand ( n3366, n26, n90 );
and ( n3367, n68, n100 );
nor ( n3368, n15, n36 );
or ( n3369, n8, n61 );
and ( n3370, n12, n140 );
or ( n3371, n21, n121 );
xor ( n3372, n74, n93 );
nor ( n3373, n0, n53 );
xor ( n3374, n62, n69 );
xor ( n3375, n43, n121 );
nor ( n3376, n30, n104 );
nor ( n3377, n43, n51 );
and ( n3378, n17, n117 );
or ( n3379, n0, n75 );
and ( n3380, n24, n86 );
xor ( n3381, n16, n71 );
xor ( n3382, n29, n140 );
and ( n3383, n11, n87 );
nor ( n3384, n58, n134 );
xor ( n3385, n107, n129 );
and ( n3386, n36, n103 );
nor ( n3387, n28, n98 );
nand ( n3388, n9, n48 );
or ( n3389, n11, n133 );
nand ( n3390, n31, n75 );
and ( n3391, n22, n57 );
xor ( n3392, n87, n130 );
nand ( n3393, n92, n135 );
or ( n3394, n59, n82 );
nand ( n3395, n101, n115 );
nor ( n3396, n63, n131 );
or ( n3397, n21, n108 );
nand ( n3398, n24, n59 );
nand ( n3399, n17, n100 );
and ( n3400, n24, n142 );
xor ( n3401, n6, n10 );
or ( n3402, n63, n124 );
or ( n3403, n93, n118 );
and ( n3404, n9, n119 );
nand ( n3405, n13, n50 );
and ( n3406, n22, n43 );
xor ( n3407, n52, n89 );
nand ( n3408, n19, n108 );
xor ( n3409, n103, n125 );
nand ( n3410, n87, n125 );
and ( n3411, n28, n93 );
xor ( n3412, n67, n72 );
or ( n3413, n83, n104 );
or ( n3414, n84, n111 );
xor ( n3415, n56, n72 );
xor ( n3416, n30, n57 );
nand ( n3417, n1, n33 );
or ( n3418, n27, n60 );
nor ( n3419, n77, n116 );
or ( n3420, n52, n65 );
nor ( n3421, n54, n132 );
nor ( n3422, n47, n103 );
or ( n3423, n45, n133 );
nor ( n3424, n53, n113 );
xor ( n3425, n5, n97 );
nand ( n3426, n16, n117 );
nand ( n3427, n60, n92 );
or ( n3428, n86, n93 );
and ( n3429, n15, n86 );
nand ( n3430, n100, n137 );
and ( n3431, n84, n90 );
xor ( n3432, n59, n99 );
xor ( n3433, n64, n95 );
xor ( n3434, n75, n135 );
nor ( n3435, n22, n110 );
nand ( n3436, n35, n90 );
nand ( n3437, n89, n101 );
nor ( n3438, n3, n20 );
xor ( n3439, n129, n132 );
or ( n3440, n52, n128 );
or ( n3441, n19, n65 );
or ( n3442, n19, n142 );
nand ( n3443, n37, n58 );
and ( n3444, n18, n78 );
nand ( n3445, n31, n67 );
nor ( n3446, n29, n45 );
xor ( n3447, n88, n119 );
nor ( n3448, n86, n137 );
and ( n3449, n28, n125 );
nor ( n3450, n75, n103 );
and ( n3451, n26, n84 );
nand ( n3452, n9, n37 );
xor ( n3453, n116, n136 );
or ( n3454, n30, n142 );
and ( n3455, n42, n82 );
nor ( n3456, n14, n117 );
xor ( n3457, n67, n73 );
nand ( n3458, n67, n96 );
nand ( n3459, n6, n59 );
or ( n3460, n106, n128 );
nor ( n3461, n10, n64 );
nand ( n3462, n38, n98 );
xor ( n3463, n59, n107 );
nand ( n3464, n5, n116 );
xor ( n3465, n29, n81 );
and ( n3466, n25, n78 );
and ( n3467, n106, n117 );
xor ( n3468, n40, n113 );
and ( n3469, n6, n138 );
nand ( n3470, n20, n44 );
and ( n3471, n48, n106 );
and ( n3472, n1, n140 );
xor ( n3473, n60, n66 );
and ( n3474, n23, n121 );
nand ( n3475, n67, n88 );
xor ( n3476, n54, n85 );
nand ( n3477, n76, n90 );
xor ( n3478, n59, n67 );
and ( n3479, n11, n88 );
nor ( n3480, n33, n87 );
nand ( n3481, n48, n140 );
nand ( n3482, n12, n73 );
or ( n3483, n9, n137 );
and ( n3484, n1, n63 );
or ( n3485, n11, n21 );
nand ( n3486, n113, n131 );
and ( n3487, n50, n108 );
or ( n3488, n82, n121 );
nor ( n3489, n30, n135 );
nand ( n3490, n62, n89 );
xor ( n3491, n0, n77 );
nand ( n3492, n38, n87 );
xor ( n3493, n12, n29 );
nor ( n3494, n41, n138 );
or ( n3495, n70, n106 );
nand ( n3496, n26, n77 );
and ( n3497, n51, n101 );
or ( n3498, n38, n131 );
nand ( n3499, n52, n86 );
xor ( n3500, n33, n119 );
and ( n3501, n50, n80 );
or ( n3502, n24, n57 );
xor ( n3503, n120, n124 );
nand ( n3504, n50, n70 );
and ( n3505, n83, n127 );
and ( n3506, n41, n95 );
nand ( n3507, n100, n105 );
nand ( n3508, n99, n124 );
or ( n3509, n86, n114 );
or ( n3510, n57, n138 );
nand ( n3511, n12, n80 );
xor ( n3512, n65, n88 );
nand ( n3513, n103, n124 );
or ( n3514, n84, n142 );
or ( n3515, n63, n68 );
and ( n3516, n16, n23 );
and ( n3517, n113, n125 );
and ( n3518, n1, n88 );
or ( n3519, n95, n105 );
and ( n3520, n45, n67 );
and ( n3521, n14, n51 );
xor ( n3522, n52, n143 );
nor ( n3523, n134, n143 );
or ( n3524, n122, n133 );
nor ( n3525, n39, n74 );
or ( n3526, n55, n112 );
xor ( n3527, n57, n127 );
xor ( n3528, n89, n106 );
or ( n3529, n80, n126 );
nand ( n3530, n20, n87 );
xor ( n3531, n21, n59 );
or ( n3532, n17, n70 );
nor ( n3533, n19, n56 );
or ( n3534, n36, n86 );
nand ( n3535, n27, n34 );
and ( n3536, n75, n138 );
nor ( n3537, n20, n139 );
xor ( n3538, n83, n128 );
nand ( n3539, n79, n97 );
xor ( n3540, n1, n35 );
nor ( n3541, n93, n95 );
xor ( n3542, n74, n85 );
or ( n3543, n35, n102 );
xor ( n3544, n57, n126 );
or ( n3545, n72, n122 );
nor ( n3546, n102, n138 );
nand ( n3547, n75, n108 );
and ( n3548, n11, n142 );
or ( n3549, n81, n82 );
or ( n3550, n4, n74 );
xor ( n3551, n109, n118 );
or ( n3552, n93, n141 );
xor ( n3553, n29, n74 );
nand ( n3554, n94, n117 );
xor ( n3555, n48, n62 );
xor ( n3556, n18, n72 );
xor ( n3557, n1, n13 );
and ( n3558, n86, n107 );
and ( n3559, n11, n39 );
nand ( n3560, n68, n98 );
xor ( n3561, n83, n143 );
nor ( n3562, n110, n122 );
and ( n3563, n122, n130 );
xor ( n3564, n30, n95 );
nor ( n3565, n77, n86 );
or ( n3566, n47, n63 );
xor ( n3567, n28, n50 );
or ( n3568, n79, n92 );
and ( n3569, n58, n124 );
xor ( n3570, n52, n76 );
nand ( n3571, n15, n38 );
nand ( n3572, n43, n123 );
nor ( n3573, n7, n93 );
or ( n3574, n13, n74 );
and ( n3575, n16, n32 );
xor ( n3576, n13, n111 );
nor ( a, n3313, n440 );
or ( b, n1565, n2293 );
nand ( c, n2785, n3368 );
nand ( d, n2938, n2017 );
xor ( e, n706, n2426 );
or ( f, n273, n152 );

not ( w1 , c );
and ( w2 , a , w1 );
nor ( w3 , a , b );
and ( w4 , b , c );
and ( w5 , c , d );
and ( y1 , b , w2 , w5);
or ( y2 , w2 , w3 , w4 );

endmodule
