module top ( in0,  in1,  in2,  in3,  in4,  in5,  in6,  in7,  in8,  in9,  in10,  in11,  in12,  in13,  in14,  in15,  in16,  in17,  in18,  in19 , i0,  i1,  i2,  i3,  i4,  i5,  i6,  i7,  i8,  i9,  i10,  i11,  i12,  i13,  i14,  i15,  i16,  i17,  i18,  i19, g11 , g12 , g13 , g14 , g15 , g16 );
input in0,  in1,  in2,  in3,  in4,  in5,  in6,  in7,  in8,  in9,  in10,  in11,  in12,  in13,  in14,  in15,  in16,  in17,  in18,  in19;
input i0,  i1,  i2,  i3,  i4,  i5,  i6,  i7,  i8,  i9,  i10,  i11,  i12,  i13,  i14,  i15,  i16,  i17,  i18,  i19;

wire g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10;
output g11 , g12 , g13 , g14 , g15 , g16 ;
wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 ,
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 ,
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 ,
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 ,
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 ,
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 ,
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 ,
     n70 , n71 , n72 , n73 ;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850;

or ( w0, in5, in17 );
or ( w1, in4, in17 );
and ( w2, in4, in18 );
nand ( w3, in2, in13 );
or ( w4, in11, in15 );
nor ( w5, in8, in13 );
and ( w6, in6, in7 );
nand ( w7, in11, in13 );
or ( w8, in8, in12 );
or ( w9, in1, in5 );
or ( w10, in0, in7 );
or ( w11, in13, in14 );
xor ( w12, in9, in11 );
or ( w13, in6, in9 );
xor ( w14, in4, in11 );
and ( w15, in8, in11 );
or ( w16, in10, in19 );
xor ( w17, in11, in19 );
or ( w18, in7, in17 );
xor ( w19, in7, in18 );
xor ( w20, in15, in16 );
xor ( w21, in0, in16 );
nand ( w22, in8, in15 );
nor ( w23, in3, in5 );
xor ( w24, in0, in5 );
and ( w25, in12, in15 );
or ( w26, in5, in10 );
or ( w27, in1, in14 );
or ( w28, in12, in14 );
nand ( w29, in4, in5 );
nand ( w30, in0, in15 );
or ( w31, in2, in14 );
nand ( w32, in8, in18 );
and ( w33, in3, in18 );
nand ( w34, in1, in15 );
and ( w35, in7, in14 );
and ( w36, in9, in12 );
nor ( w37, in7, in19 );
nor ( w38, in0, in4 );
xor ( w39, in10, in17 );
nand ( w40, in7, in11 );
and ( w41, in4, in15 );
nand ( w42, in0, in19 );
nand ( w43, in3, in10 );
and ( w44, in12, in16 );
or ( w45, in12, in17 );
nor ( w46, in16, in17 );
or ( w47, in2, in18 );
and ( w48, in6, in10 );
nand ( w49, in9, in15 );
and ( w50, in1, in8 );
and ( w51, in9, in14 );
and ( w52, in16, in19 );
nand ( w53, in2, in12 );
or ( w54, in9, in13 );
and ( w55, in14, in15 );
or ( w56, in4, in9 );
and ( w57, in8, in17 );
xor ( w58, in1, in16 );
or ( w59, in2, in15 );
xor ( w60, in6, in15 );
nand ( w61, in0, in2 );
nand ( w62, in0, in12 );
or ( w63, w31, w50 );
or ( w64, w14, w48 );
nand ( w65, w13, w42 );
nor ( w66, w33, w49 );
nor ( w67, w33, w46 );
or ( w68, w34, w60 );
nand ( w69, w23, w42 );
xor ( w70, w11, w16 );
nor ( w71, w15, w16 );
or ( w72, w16, w18 );
nor ( w73, w11, w23 );
xor ( w74, w30, w54 );
nor ( w75, w9, w41 );
and ( w76, w4, w36 );
xor ( w77, w24, w33 );
nor ( w78, w5, w49 );
xor ( w79, w51, w58 );
xor ( w80, w53, w57 );
or ( w81, w31, w46 );
or ( w82, w34, w61 );
xor ( w83, w10, w47 );
and ( w84, w8, w60 );
nand ( w85, w45, w53 );
or ( w86, w30, w58 );
and ( w87, w3, w5 );
and ( w88, w2, w46 );
or ( w89, w19, w50 );
and ( w90, w1, w10 );
nor ( w91, w3, w53 );
and ( w92, w19, w26 );
xor ( w93, w2, w28 );
nor ( w94, w7, w14 );
xor ( w95, w3, w14 );
nor ( w96, w18, w31 );
and ( w97, w7, w44 );
xor ( w98, w23, w29 );
nand ( w99, w13, w31 );
nand ( w100, w24, w60 );
xor ( w101, w16, w17 );
or ( w102, w34, w51 );
and ( w103, w15, w25 );
and ( w104, w18, w28 );
nand ( w105, w5, w25 );
nor ( w106, w18, w21 );
or ( w107, w38, w76 );
or ( w108, w3, w56 );
nor ( w109, w39, w47 );
and ( w110, w67, w75 );
nand ( w111, w0, w38 );
nor ( w112, w1, w37 );
nand ( w113, w66, w86 );
and ( w114, w30, w63 );
and ( w115, w7, w91 );
and ( w116, w29, w64 );
or ( w117, w10, w24 );
nor ( w118, w27, w90 );
or ( w119, w68, w92 );
and ( w120, w6, w8 );
nand ( w121, w43, w67 );
nor ( w122, w37, w72 );
and ( w123, w60, w79 );
xor ( w124, w12, w29 );
or ( w125, w22, w39 );
nand ( w126, w54, w76 );
or ( w127, w69, w71 );
and ( w128, w8, w84 );
and ( w129, w28, w99 );
or ( w130, w24, w91 );
nor ( w131, w65, w79 );
and ( w132, w55, w78 );
nor ( w133, w101, w103 );
or ( w134, w75, w90 );
xor ( w135, w30, w39 );
xor ( w136, w0, w8 );
nor ( w137, w35, w48 );
or ( w138, w28, w74 );
and ( w139, w18, w85 );
nand ( w140, w95, w98 );
or ( w141, w82, w90 );
xor ( w142, w59, w68 );
and ( w143, w25, w88 );
and ( w144, w15, w55 );
nand ( w145, w10, w17 );
and ( w146, w61, w96 );
xor ( w147, w30, w102 );
or ( w148, w37, w43 );
xor ( w149, w71, w102 );
and ( w150, w30, w31 );
xor ( w151, w33, w59 );
or ( w152, w73, w94 );
nand ( w153, w0, w99 );
xor ( w154, w58, w88 );
and ( w155, w91, w92 );
and ( w156, w38, w56 );
nand ( w157, w24, w61 );
or ( w158, w41, w62 );
or ( w159, w39, w103 );
xor ( w160, w25, w95 );
xor ( w161, w31, w33 );
and ( w162, w74, w92 );
nor ( w163, w3, w86 );
or ( w164, w50, w55 );
nand ( w165, w33, w98 );
or ( w166, w26, w33 );
or ( w167, w35, w81 );
or ( w168, w30, w83 );
or ( w169, w56, w61 );
nor ( w170, w8, w13 );
nand ( w171, w25, w30 );
nor ( w172, w32, w75 );
nand ( w173, w21, w89 );
xor ( w174, w53, w67 );
xor ( w175, w27, w44 );
nor ( w176, w57, w159 );
and ( w177, w59, w125 );
or ( w178, w43, w70 );
nor ( w179, w32, w147 );
xor ( w180, w132, w169 );
or ( w181, w51, w91 );
nand ( w182, w63, w146 );
xor ( w183, w39, w138 );
xor ( w184, w52, w134 );
and ( w185, w49, w124 );
nand ( w186, w29, w104 );
nor ( w187, w89, w131 );
or ( w188, w80, w121 );
and ( w189, w66, w140 );
and ( w190, w26, w134 );
nor ( w191, w72, w90 );
xor ( w192, w75, w91 );
or ( w193, w27, w34 );
or ( w194, w134, w147 );
nor ( w195, w5, w163 );
or ( w196, w108, w163 );
and ( w197, w27, w98 );
nand ( w198, w110, w137 );
nand ( w199, w17, w165 );
or ( w200, w5, w142 );
nor ( w201, w5, w119 );
and ( w202, w13, w162 );
xor ( w203, w81, w110 );
nand ( w204, w154, w171 );
nand ( w205, w6, w37 );
nand ( w206, w52, w119 );
nor ( w207, w6, w67 );
or ( w208, w71, w72 );
and ( w209, w63, w65 );
nand ( w210, w41, w111 );
or ( w211, w57, w142 );
or ( w212, w59, w74 );
nor ( w213, w77, w162 );
and ( w214, w15, w110 );
or ( w215, w88, w149 );
and ( w216, w7, w38 );
nor ( w217, w20, w42 );
nor ( w218, w9, w26 );
xor ( w219, w9, w160 );
nor ( w220, w56, w107 );
or ( w221, w25, w136 );
xor ( w222, w47, w82 );
or ( w223, w89, w116 );
or ( w224, w91, w170 );
xor ( w225, w30, w101 );
nor ( w226, w67, w130 );
or ( w227, w33, w37 );
and ( w228, w72, w118 );
and ( w229, w75, w76 );
nand ( w230, w98, w173 );
nand ( w231, w98, w166 );
and ( w232, w91, w103 );
nor ( w233, w65, w124 );
xor ( w234, w15, w117 );
nor ( w235, w0, w162 );
or ( w236, w45, w95 );
and ( w237, w19, w123 );
nand ( w238, w15, w165 );
nand ( w239, w19, w91 );
nor ( w240, w66, w134 );
nor ( w241, w5, w127 );
nor ( w242, w15, w101 );
nor ( w243, w66, w89 );
nor ( w244, w137, w164 );
nor ( w245, w136, w174 );
nand ( w246, w35, w101 );
and ( w247, w20, w35 );
and ( w248, w69, w97 );
xor ( w249, w150, w167 );
or ( w250, w65, w132 );
nand ( w251, w60, w81 );
xor ( w252, w35, w105 );
nor ( w253, w131, w132 );
nand ( w254, w9, w118 );
and ( w255, w60, w169 );
or ( w256, w20, w87 );
nand ( w257, w20, w122 );
nand ( w258, w43, w167 );
xor ( w259, w8, w124 );
nor ( w260, w115, w126 );
nor ( w261, w0, w119 );
xor ( w262, w7, w118 );
or ( w263, w90, w119 );
nor ( w264, w32, w166 );
nor ( w265, w76, w169 );
xor ( w266, w37, w123 );
nand ( w267, w22, w145 );
xor ( w268, w156, w173 );
nand ( w269, w75, w113 );
or ( w270, w34, w90 );
nor ( w271, w95, w115 );
or ( w272, w20, w79 );
and ( w273, w110, w131 );
nor ( w274, w119, w153 );
nor ( w275, w32, w109 );
and ( w276, w38, w109 );
xor ( w277, w31, w79 );
xor ( w278, w86, w104 );
nor ( w279, w31, w137 );
xor ( w280, w58, w119 );
nor ( w281, w62, w70 );
xor ( w282, w86, w110 );
or ( w283, w19, w83 );
and ( w284, w99, w100 );
or ( w285, w28, w87 );
or ( w286, w101, w108 );
and ( w287, w134, w151 );
xor ( w288, w115, w132 );
or ( w289, w128, w170 );
and ( w290, w40, w129 );
nor ( w291, w38, w144 );
or ( w292, w0, w48 );
nand ( w293, w60, w74 );
nand ( w294, w127, w174 );
and ( w295, w137, w172 );
xor ( w296, w2, w48 );
nand ( w297, w176, w199 );
nor ( w298, w6, w24 );
and ( w299, w125, w215 );
and ( w300, w72, w272 );
or ( w301, w197, w288 );
and ( w302, w7, w88 );
and ( w303, w110, w217 );
nor ( w304, w23, w115 );
nand ( w305, w157, w225 );
or ( w306, w164, w228 );
or ( w307, w219, w264 );
and ( w308, w63, w190 );
and ( w309, w196, w232 );
xor ( w310, w229, w266 );
or ( w311, w5, w228 );
or ( w312, w195, w256 );
nand ( w313, w181, w292 );
or ( w314, w135, w266 );
and ( w315, w170, w255 );
or ( w316, w37, w126 );
nor ( w317, w286, w291 );
xor ( w318, w43, w212 );
and ( w319, w72, w273 );
or ( w320, w35, w263 );
nor ( w321, w85, w259 );
nand ( w322, w70, w103 );
and ( w323, w198, w235 );
xor ( w324, w3, w174 );
or ( w325, w185, w274 );
or ( w326, w17, w121 );
xor ( w327, w102, w122 );
and ( w328, w138, w227 );
or ( w329, w16, w26 );
xor ( w330, w124, w187 );
nand ( w331, w117, w124 );
xor ( w332, w94, w186 );
nand ( w333, w233, w244 );
or ( w334, w143, w253 );
nor ( w335, w113, w119 );
xor ( w336, w204, w282 );
xor ( w337, w6, w141 );
nor ( w338, w157, w248 );
and ( w339, w177, w295 );
or ( w340, w255, w294 );
nand ( w341, w0, w284 );
xor ( w342, w85, w105 );
and ( w343, w108, w147 );
nand ( w344, w39, w83 );
or ( w345, w82, w295 );
and ( w346, w12, w103 );
nor ( w347, w68, w79 );
or ( w348, w0, w186 );
or ( w349, w206, w280 );
nor ( w350, w129, w157 );
and ( w351, w159, w289 );
nor ( w352, w31, w292 );
xor ( w353, w145, w278 );
or ( w354, w150, w177 );
or ( w355, w150, w288 );
and ( w356, w69, w262 );
xor ( w357, w231, w252 );
xor ( w358, w126, w139 );
nand ( w359, w82, w240 );
nor ( w360, w33, w144 );
and ( w361, w117, w143 );
and ( w362, w50, w85 );
nand ( w363, w173, w177 );
nand ( w364, w73, w243 );
xor ( w365, w1, w88 );
nor ( w366, w120, w148 );
nand ( w367, w67, w95 );
nand ( w368, w202, w221 );
and ( w369, w232, w235 );
xor ( w370, w114, w126 );
xor ( w371, w31, w250 );
xor ( w372, w26, w242 );
or ( w373, w47, w231 );
xor ( w374, w245, w251 );
or ( w375, w219, w283 );
xor ( w376, w121, w230 );
nor ( w377, w28, w153 );
xor ( w378, w30, w98 );
and ( w379, w109, w265 );
xor ( w380, w248, w269 );
nor ( w381, w77, w134 );
xor ( w382, w204, w254 );
xor ( w383, w125, w242 );
and ( w384, w123, w263 );
xor ( w385, w198, w274 );
nor ( w386, w113, w282 );
nor ( w387, w46, w108 );
and ( w388, w88, w207 );
and ( w389, w83, w88 );
or ( w390, w170, w176 );
or ( w391, w42, w254 );
nand ( w392, w187, w272 );
and ( w393, w135, w160 );
nor ( w394, w127, w282 );
and ( w395, w40, w58 );
and ( w396, w167, w228 );
nand ( w397, w89, w190 );
and ( w398, w63, w200 );
or ( w399, w74, w212 );
nand ( w400, w252, w274 );
and ( w401, w47, w166 );
xor ( w402, w191, w260 );
or ( w403, w101, w217 );
nand ( w404, w24, w36 );
or ( w405, w245, w292 );
xor ( w406, w45, w209 );
and ( w407, w60, w294 );
and ( w408, w32, w214 );
or ( w409, w73, w229 );
and ( w410, w7, w26 );
nand ( w411, w164, w210 );
xor ( w412, w23, w173 );
xor ( w413, w74, w257 );
nand ( w414, w107, w294 );
nand ( w415, w67, w202 );
xor ( w416, w154, w180 );
xor ( w417, w156, w207 );
or ( w418, w149, w236 );
and ( w419, w133, w288 );
nor ( w420, w20, w205 );
xor ( w421, w9, w172 );
xor ( w422, w276, w289 );
nand ( w423, w9, w217 );
and ( w424, w61, w90 );
or ( w425, w101, w132 );
nand ( w426, w112, w277 );
or ( w427, w48, w98 );
nand ( w428, w182, w249 );
nor ( w429, w4, w7 );
xor ( w430, w113, w139 );
nand ( w431, w21, w152 );
or ( w432, w76, w234 );
xor ( w433, w139, w170 );
and ( w434, w121, w277 );
or ( w435, w130, w290 );
nor ( w436, w139, w171 );
and ( w437, w81, w127 );
and ( w438, w6, w98 );
and ( w439, w36, w192 );
nand ( w440, w75, w242 );
or ( w441, w194, w273 );
xor ( w442, w122, w287 );
xor ( w443, w151, w233 );
nor ( w444, w193, w234 );
nor ( w445, w157, w217 );
nand ( w446, w32, w58 );
nand ( w447, w219, w252 );
or ( w448, w4, w205 );
and ( w449, w49, w230 );
xor ( w450, w114, w221 );
or ( w451, w75, w101 );
xor ( w452, w8, w265 );
or ( w453, w160, w284 );
and ( w454, w197, w200 );
or ( w455, w178, w185 );
nor ( w456, w74, w190 );
nand ( w457, w150, w170 );
and ( w458, w37, w262 );
or ( w459, w138, w148 );
and ( w460, w66, w99 );
nor ( w461, w31, w258 );
and ( w462, w147, w241 );
nor ( w463, w1, w65 );
nand ( w464, w54, w277 );
nand ( w465, w62, w91 );
nor ( w466, w165, w224 );
nand ( w467, w108, w197 );
or ( w468, w46, w138 );
and ( w469, w35, w112 );
xor ( w470, w50, w205 );
nand ( w471, w281, w290 );
nand ( w472, w49, w75 );
or ( w473, w3, w98 );
and ( w474, w15, w41 );
nand ( w475, w28, w269 );
and ( w476, w23, w201 );
and ( w477, w95, w195 );
and ( w478, w40, w230 );
or ( w479, w20, w146 );
xor ( w480, w61, w146 );
nor ( w481, w61, w261 );
nand ( w482, w87, w261 );
xor ( w483, w162, w274 );
nor ( w484, w40, w134 );
xor ( w485, w230, w289 );
nor ( w486, w276, w282 );
xor ( w487, w83, w262 );
and ( w488, w247, w262 );
and ( w489, w111, w152 );
nand ( w490, w197, w254 );
nand ( w491, w176, w180 );
or ( w492, w93, w186 );
nand ( w493, w45, w245 );
nor ( w494, w202, w280 );
nor ( w495, w161, w180 );
nand ( w496, w179, w280 );
nand ( w497, w16, w214 );
nor ( w498, w44, w98 );
and ( w499, w2, w217 );
nand ( w500, w53, w109 );
or ( w501, w70, w144 );
and ( w502, w93, w489 );
xor ( w503, w107, w159 );
nor ( w504, w323, w435 );
xor ( w505, w282, w480 );
or ( w506, w183, w196 );
and ( w507, w13, w47 );
and ( w508, w415, w471 );
xor ( w509, w265, w410 );
xor ( w510, w82, w218 );
or ( w511, w69, w314 );
or ( w512, w90, w111 );
nand ( w513, w30, w444 );
nand ( w514, w438, w452 );
or ( w515, w246, w394 );
or ( w516, w370, w496 );
xor ( w517, w196, w496 );
or ( w518, w113, w481 );
or ( w519, w7, w449 );
and ( w520, w403, w464 );
xor ( w521, w22, w310 );
and ( w522, w334, w461 );
xor ( w523, w179, w272 );
nand ( w524, w262, w375 );
and ( w525, w8, w299 );
nor ( w526, w366, w468 );
nand ( w527, w217, w481 );
xor ( w528, w11, w235 );
nor ( w529, w206, w403 );
nand ( w530, w126, w360 );
and ( w531, w85, w467 );
xor ( w532, w9, w64 );
xor ( w533, w291, w436 );
and ( w534, w26, w148 );
and ( w535, w345, w458 );
or ( w536, w123, w187 );
nand ( w537, w29, w105 );
nand ( w538, w85, w421 );
nand ( w539, w141, w439 );
and ( w540, w218, w245 );
nor ( w541, w19, w362 );
nand ( w542, w51, w177 );
nand ( w543, w105, w341 );
and ( w544, w305, w387 );
and ( w545, w248, w325 );
xor ( w546, w103, w151 );
nand ( w547, w42, w409 );
or ( w548, w48, w75 );
and ( w549, w121, w220 );
xor ( w550, w236, w331 );
or ( w551, w334, w483 );
xor ( w552, w59, w294 );
or ( w553, w368, w395 );
or ( w554, w277, w445 );
nor ( w555, w136, w268 );
and ( w556, w256, w390 );
nor ( w557, w103, w467 );
xor ( w558, w128, w444 );
or ( w559, w227, w373 );
or ( w560, w47, w122 );
and ( w561, w133, w281 );
and ( w562, w50, w297 );
nand ( w563, w128, w429 );
nand ( w564, w266, w497 );
and ( w565, w304, w342 );
nor ( w566, w204, w339 );
or ( w567, w318, w441 );
nor ( w568, w91, w346 );
or ( w569, w44, w192 );
and ( w570, w151, w443 );
or ( w571, w178, w184 );
and ( w572, w437, w470 );
and ( w573, w116, w349 );
and ( w574, w12, w372 );
nand ( w575, w174, w458 );
xor ( w576, w204, w250 );
nor ( w577, w258, w365 );
and ( w578, w133, w427 );
nor ( w579, w76, w119 );
xor ( w580, w19, w22 );
xor ( w581, w469, w493 );
nor ( w582, w159, w337 );
nand ( w583, w136, w254 );
and ( w584, w90, w489 );
xor ( w585, w113, w247 );
nand ( w586, w183, w252 );
and ( w587, w89, w308 );
or ( w588, w28, w459 );
and ( w589, w15, w376 );
nand ( w590, w273, w316 );
nand ( w591, w265, w316 );
and ( w592, w182, w425 );
xor ( w593, w340, w497 );
xor ( w594, w182, w372 );
and ( w595, w125, w197 );
nor ( w596, w150, w382 );
nand ( w597, w413, w459 );
or ( w598, w215, w397 );
xor ( w599, w3, w121 );
and ( w600, w17, w146 );
nand ( w601, w111, w199 );
or ( w602, w277, w412 );
nand ( w603, w196, w218 );
nand ( w604, w352, w460 );
nand ( w605, w39, w346 );
nor ( w606, w341, w387 );
or ( w607, w53, w454 );
nand ( w608, w239, w417 );
or ( w609, w26, w69 );
nand ( w610, w336, w387 );
or ( w611, w15, w426 );
and ( w612, w85, w126 );
and ( w613, w286, w447 );
nor ( w614, w83, w485 );
nand ( w615, w196, w427 );
nor ( w616, w141, w187 );
nand ( w617, w174, w448 );
nand ( w618, w352, w355 );
or ( w619, w111, w273 );
nor ( w620, w360, w402 );
and ( w621, w279, w380 );
xor ( w622, w267, w463 );
nand ( w623, w214, w277 );
nor ( w624, w87, w254 );
nand ( w625, w108, w367 );
or ( w626, w211, w392 );
nand ( w627, w27, w131 );
nand ( w628, w68, w385 );
or ( w629, w73, w279 );
nand ( w630, w99, w471 );
or ( w631, w383, w492 );
nand ( w632, w222, w468 );
and ( w633, w109, w469 );
xor ( w634, w346, w485 );
nand ( w635, w8, w185 );
or ( w636, w286, w319 );
and ( w637, w446, w482 );
or ( w638, w347, w466 );
nand ( w639, w218, w345 );
nand ( w640, w224, w471 );
and ( w641, w192, w335 );
and ( w642, w270, w279 );
nand ( w643, w71, w137 );
nor ( w644, w107, w163 );
xor ( w645, w73, w499 );
xor ( w646, w49, w434 );
or ( w647, w39, w285 );
or ( w648, w91, w93 );
nand ( w649, w14, w207 );
xor ( w650, w132, w468 );
nand ( w651, w318, w444 );
xor ( w652, w269, w441 );
and ( w653, w45, w93 );
xor ( w654, w58, w497 );
xor ( w655, w150, w454 );
or ( w656, w67, w173 );
or ( w657, w331, w417 );
nor ( w658, w159, w489 );
nor ( w659, w147, w327 );
or ( w660, w306, w460 );
nand ( w661, w383, w477 );
and ( w662, w409, w464 );
xor ( w663, w285, w394 );
xor ( w664, w275, w367 );
and ( w665, w385, w488 );
and ( w666, w413, w488 );
or ( w667, w72, w87 );
nand ( w668, w260, w443 );
and ( w669, w128, w176 );
xor ( w670, w340, w448 );
nand ( w671, w395, w475 );
or ( w672, w214, w482 );
xor ( w673, w85, w339 );
and ( w674, w401, w448 );
xor ( w675, w179, w387 );
or ( w676, w33, w313 );
nor ( w677, w233, w465 );
or ( w678, w125, w163 );
nor ( w679, w250, w362 );
xor ( w680, w10, w173 );
or ( w681, w190, w404 );
nand ( w682, w50, w319 );
nand ( w683, w262, w313 );
xor ( w684, w488, w500 );
and ( w685, w120, w441 );
nor ( w686, w124, w162 );
or ( w687, w232, w409 );
nand ( w688, w3, w350 );
or ( w689, w48, w368 );
nand ( w690, w382, w500 );
or ( w691, w72, w352 );
xor ( w692, w52, w119 );
nand ( w693, w177, w251 );
nor ( w694, w45, w347 );
and ( w695, w7, w18 );
xor ( w696, w365, w446 );
nor ( w697, w58, w96 );
or ( w698, w61, w146 );
and ( w699, w45, w179 );
and ( w700, w252, w476 );
nand ( w701, w65, w448 );
or ( w702, w175, w378 );
and ( w703, w225, w348 );
xor ( w704, w7, w495 );
or ( w705, w63, w402 );
xor ( w706, w33, w198 );
nor ( w707, w397, w437 );
xor ( w708, w352, w408 );
and ( w709, w134, w309 );
and ( w710, w77, w237 );
and ( w711, w254, w383 );
nand ( w712, w150, w497 );
nand ( w713, w411, w461 );
and ( w714, w100, w359 );
and ( w715, w91, w235 );
xor ( w716, w110, w442 );
xor ( w717, w130, w258 );
and ( w718, w204, w270 );
nor ( w719, w383, w467 );
nand ( w720, w266, w499 );
or ( w721, w231, w319 );
or ( w722, w161, w323 );
or ( w723, w102, w415 );
xor ( w724, w79, w405 );
nor ( w725, w370, w451 );
and ( w726, w25, w55 );
and ( w727, w313, w414 );
and ( w728, w30, w263 );
and ( w729, w122, w293 );
xor ( w730, w272, w305 );
nand ( w731, w69, w442 );
or ( w732, w15, w454 );
and ( w733, w224, w273 );
nor ( w734, w460, w465 );
xor ( w735, w365, w433 );
xor ( w736, w50, w374 );
xor ( w737, w223, w408 );
xor ( w738, w64, w274 );
or ( w739, w89, w390 );
nand ( w740, w400, w479 );
nand ( w741, w339, w340 );
and ( w742, w75, w364 );
or ( w743, w79, w469 );
and ( w744, w166, w204 );
and ( w745, w386, w476 );
xor ( w746, w54, w180 );
nor ( w747, w296, w374 );
xor ( w748, w420, w467 );
or ( w749, w34, w461 );
xor ( w750, w60, w279 );
nand ( w751, w128, w432 );
and ( w752, w41, w333 );
or ( w753, w192, w375 );
or ( w754, w231, w498 );
and ( w755, w336, w456 );
nor ( w756, w28, w220 );
and ( w757, w219, w269 );
nand ( w758, w126, w172 );
and ( w759, w34, w39 );
and ( w760, w322, w422 );
and ( w761, w179, w400 );
xor ( w762, w169, w368 );
xor ( w763, w192, w340 );
nand ( w764, w55, w64 );
nand ( w765, w16, w433 );
or ( w766, w31, w243 );
nor ( w767, w296, w426 );
xor ( w768, w348, w376 );
nor ( w769, w60, w265 );
nor ( w770, w268, w496 );
and ( w771, w208, w379 );
or ( w772, w253, w380 );
nor ( w773, w107, w329 );
nand ( w774, w322, w348 );
xor ( w775, w100, w392 );
nand ( w776, w127, w288 );
nor ( w777, w244, w409 );
nor ( w778, w107, w283 );
or ( w779, w174, w233 );
nor ( w780, w151, w276 );
or ( w781, w242, w452 );
and ( w782, w98, w418 );
nor ( w783, w82, w388 );
xor ( w784, w357, w493 );
and ( w785, w238, w491 );
xor ( w786, w178, w313 );
nand ( w787, w114, w301 );
nor ( w788, w216, w277 );
nor ( w789, w169, w203 );
xor ( w790, w42, w54 );
and ( w791, w413, w465 );
xor ( w792, w83, w215 );
and ( w793, w183, w469 );
nand ( w794, w408, w432 );
or ( w795, w290, w320 );
and ( w796, w49, w466 );
xor ( w797, w122, w310 );
nor ( w798, w61, w432 );
nor ( w799, w422, w446 );
xor ( w800, w19, w264 );
and ( w801, w164, w434 );
or ( w802, w336, w492 );
and ( w803, w270, w370 );
nand ( w804, w292, w411 );
or ( w805, w47, w345 );
nand ( w806, w322, w324 );
and ( w807, w53, w81 );
nor ( w808, w328, w379 );
nor ( w809, w360, w480 );
nor ( w810, w94, w121 );
xor ( w811, w45, w327 );
nor ( w812, w52, w402 );
nor ( w813, w115, w262 );
nor ( w814, w241, w484 );
or ( w815, w335, w337 );
nand ( w816, w164, w303 );
and ( w817, w398, w430 );
xor ( w818, w21, w173 );
or ( w819, w331, w395 );
nor ( w820, w187, w288 );
and ( w821, w101, w249 );
or ( w822, w259, w325 );
nor ( w823, w121, w486 );
or ( w824, w332, w446 );
nand ( w825, w115, w319 );
and ( w826, w260, w486 );
nand ( w827, w169, w217 );
xor ( w828, w173, w255 );
and ( w829, w26, w90 );
or ( w830, w87, w451 );
and ( w831, w64, w303 );
nor ( w832, w25, w433 );
nor ( w833, w121, w162 );
or ( w834, w84, w388 );
nor ( w835, w98, w487 );
nor ( w836, w401, w461 );
nand ( w837, w86, w208 );
nand ( w838, w32, w286 );
nand ( w839, w256, w366 );
xor ( w840, w93, w168 );
xor ( w841, w199, w203 );
nor ( w842, w50, w343 );
xor ( w843, w13, w240 );
or ( w844, w61, w350 );
and ( w845, w143, w493 );
nor ( w846, w406, w435 );
nand ( w847, w29, w138 );
or ( w848, w354, w372 );
or ( w849, w282, w348 );
xor ( w850, w115, w410 );
or ( g0, w542, w807 );
or ( g1, w605, w697 );
nor ( g2, w701, w734 );
nand ( g3, w678, w677 );
nand ( g4, w836, w821 );
or ( g5, w810, w665 );
nand ( g6, w505, w542 );
xor ( g7, w810, w550 );
and ( g8, w634, w580 );
nand ( g9, w707, w611 );
and ( g10, w668, w562 );

buf ( n1  , g0 );
buf ( n2  , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( g11 , n12  );
buf ( g12 , n13  );
buf ( g13 , n14  );
buf ( g14 , n15  );
buf ( g15 , n16  );
buf ( g16 , n17  );
buf ( n12 , n44 );
buf ( n13 , n57 );
buf ( n14 , n73 );
buf ( n15 , n50 );
buf ( n16 , n61 );
buf ( n17 , n68 );
xor ( n20 , n2 , n6 );
not ( n21 , n20 );
nand ( n22 , n4 , n8 );
nand ( n23 , n3 , n7 );
and ( n24 , n22 , n23 );
nor ( n25 , n3 , n7 );
nor ( n26 , n24 , n25 );
not ( n27 , n26 );
or ( n28 , n21 , n27 );
and ( n29 , n22 , n23 );
nor ( n30 , n29 , n25 );
or ( n31 , n20 , n30 );
nand ( n32 , n28 , n31 );
not ( n33 , n9 );
and ( n34 , n10 , n33 );
not ( n35 , n10 );
and ( n36 , n35 , n9 );
nor ( n37 , n34 , n36 );
not ( n38 , n37 );
not ( n39 , n38 );
or ( n40 , n32 , n39 );
not ( n41 , n37 );
not ( n42 , n2 );
or ( n43 , n41 , n42 );
nand ( n44 , n40 , n43 );
or ( n45 , n32 , n41 );
not ( n46 , n37 );
not ( n47 , n46 );
not ( n48 , n6 );
or ( n49 , n47 , n48 );
nand ( n50 , n45 , n49 );
xor ( n51 , n3 , n7 );
nand ( n52 , n4 , n8 );
xor ( n53 , n51 , n52 );
or ( n54 , n39 , n53 );
not ( n55 , n3 );
or ( n56 , n41 , n55 );
nand ( n57 , n54 , n56 );
or ( n58 , n53 , n41 );
not ( n59 , n7 );
or ( n60 , n47 , n59 );
nand ( n61 , n58 , n60 );
not ( n62 , n8 );
not ( n63 , n46 );
or ( n64 , n62 , n63 );
or ( n65 , n4 , n8 );
nand ( n66 , n65 , n22 );
or ( n67 , n38 , n66 );
nand ( n68 , n64 , n67 );
not ( n69 , n37 );
not ( n70 , n4 );
or ( n71 , n69 , n70 );
or ( n72 , n66 , n37 );
nand ( n73 , n71 , n72 );

wire ou0,  ou1,  ou2,  ou3,  ou4,  ou5,  ou6,  ou7,  ou8,  ou9,  ou10;
wire wi0, wi1, wi2, wi3, wi4, wi5, wi6, wi7, wi8, wi9, wi10, wi11, wi12, wi13, wi14, wi15, wi16, wi17, wi18, wi19, wi20, wi21, wi22, wi23, wi24, wi25, wi26, wi27, wi28, wi29, wi30, wi31, wi32, wi33, wi34, wi35, wi36, wi37, wi38, wi39, wi40, wi41, wi42, wi43, wi44, wi45, wi46, wi47, wi48, wi49, wi50, wi51, wi52, wi53, wi54, wi55, wi56, wi57, wi58, wi59, wi60, wi61, wi62, wi63, wi64, wi65, wi66, wi67, wi68, wi69, wi70, wi71, wi72, wi73, wi74, wi75, wi76, wi77, wi78, wi79, wi80, wi81, wi82, wi83, wi84, wi85, wi86, wi87, wi88, wi89, wi90, wi91, wi92, wi93, wi94, wi95, wi96, wi97, wi98, wi99, wi100, wi101, wi102, wi103, wi104, wi105, wi106, wi107, wi108, wi109, wi110, wi111, wi112, wi113, wi114, wi115, wi116, wi117, wi118, wi119, wi120, wi121, wi122, wi123, wi124, wi125, wi126, wi127, wi128, wi129, wi130, wi131, wi132, wi133, wi134, wi135, wi136, wi137, wi138, wi139, wi140, wi141, wi142, wi143, wi144, wi145, wi146, wi147, wi148, wi149, wi150, wi151, wi152, wi153, wi154, wi155, wi156, wi157, wi158, wi159, wi160, wi161, wi162, wi163, wi164, wi165, wi166, wi167, wi168, wi169, wi170, wi171, wi172, wi173, wi174, wi175, wi176, wi177, wi178, wi179, wi180, wi181, wi182, wi183, wi184, wi185, wi186, wi187, wi188, wi189, wi190, wi191, wi192, wi193, wi194, wi195, wi196, wi197, wi198, wi199, wi200, wi201, wi202, wi203, wi204, wi205, wi206, wi207, wi208, wi209, wi210, wi211, wi212, wi213, wi214, wi215, wi216, wi217, wi218, wi219, wi220, wi221, wi222, wi223, wi224, wi225, wi226, wi227, wi228, wi229, wi230, wi231, wi232, wi233, wi234, wi235, wi236, wi237, wi238, wi239, wi240, wi241, wi242, wi243, wi244, wi245, wi246, wi247, wi248, wi249, wi250, wi251, wi252, wi253, wi254, wi255, wi256, wi257, wi258, wi259, wi260, wi261, wi262, wi263, wi264, wi265, wi266, wi267, wi268, wi269, wi270, wi271, wi272, wi273, wi274, wi275, wi276, wi277, wi278, wi279, wi280, wi281, wi282, wi283, wi284, wi285, wi286, wi287, wi288, wi289, wi290, wi291, wi292, wi293, wi294, wi295, wi296, wi297, wi298, wi299, wi300, wi301, wi302, wi303, wi304, wi305, wi306, wi307, wi308, wi309, wi310, wi311, wi312, wi313, wi314, wi315, wi316, wi317, wi318, wi319, wi320, wi321, wi322, wi323, wi324, wi325, wi326, wi327, wi328, wi329, wi330, wi331, wi332, wi333, wi334, wi335, wi336, wi337, wi338, wi339, wi340, wi341, wi342, wi343, wi344, wi345, wi346, wi347, wi348, wi349, wi350, wi351, wi352, wi353, wi354, wi355, wi356, wi357, wi358, wi359, wi360, wi361, wi362, wi363, wi364, wi365, wi366, wi367, wi368, wi369, wi370, wi371, wi372, wi373, wi374, wi375, wi376, wi377, wi378, wi379, wi380, wi381, wi382, wi383, wi384, wi385, wi386, wi387, wi388, wi389, wi390, wi391, wi392, wi393, wi394, wi395, wi396, wi397, wi398, wi399, wi400, wi401, wi402, wi403, wi404, wi405, wi406, wi407, wi408, wi409, wi410, wi411, wi412, wi413, wi414, wi415, wi416, wi417, wi418, wi419, wi420, wi421, wi422, wi423, wi424, wi425, wi426, wi427, wi428, wi429, wi430, wi431, wi432, wi433, wi434, wi435, wi436, wi437, wi438, wi439, wi440, wi441, wi442, wi443, wi444, wi445, wi446, wi447, wi448, wi449, wi450, wi451, wi452, wi453, wi454, wi455, wi456, wi457, wi458, wi459, wi460, wi461, wi462, wi463, wi464, wi465, wi466, wi467, wi468, wi469, wi470, wi471, wi472, wi473, wi474, wi475, wi476, wi477, wi478, wi479, wi480, wi481, wi482, wi483, wi484, wi485, wi486, wi487, wi488, wi489, wi490, wi491, wi492, wi493, wi494, wi495, wi496, wi497, wi498, wi499, wi500, wi501, wi502, wi503, wi504, wi505, wi506, wi507, wi508, wi509, wi510, wi511, wi512, wi513, wi514, wi515, wi516, wi517, wi518, wi519, wi520, wi521, wi522, wi523, wi524, wi525, wi526, wi527, wi528, wi529, wi530, wi531, wi532, wi533, wi534, wi535, wi536, wi537, wi538, wi539, wi540, wi541, wi542, wi543, wi544, wi545, wi546, wi547, wi548, wi549, wi550, wi551, wi552, wi553, wi554, wi555, wi556, wi557, wi558, wi559, wi560, wi561, wi562, wi563, wi564, wi565, wi566, wi567, wi568, wi569, wi570, wi571, wi572, wi573, wi574, wi575, wi576, wi577, wi578, wi579, wi580, wi581, wi582, wi583, wi584, wi585, wi586, wi587, wi588, wi589, wi590, wi591, wi592, wi593, wi594, wi595, wi596, wi597, wi598, wi599, wi600, wi601, wi602, wi603, wi604, wi605, wi606, wi607, wi608, wi609, wi610, wi611, wi612, wi613, wi614, wi615, wi616, wi617, wi618, wi619, wi620, wi621, wi622, wi623, wi624, wi625, wi626, wi627, wi628, wi629, wi630, wi631, wi632, wi633, wi634, wi635, wi636, wi637, wi638, wi639, wi640, wi641, wi642, wi643, wi644, wi645, wi646, wi647, wi648, wi649, wi650, wi651, wi652, wi653, wi654, wi655, wi656, wi657, wi658;

and ( wi0, i4, i16 );
and ( wi1, i14, i19 );
or ( wi2, i2, i14 );
and ( wi3, i10, i17 );
and ( wi4, i7, i15 );
xor ( wi5, i8, i11 );
nand ( wi6, i7, i17 );
nor ( wi7, i9, i17 );
and ( wi8, i1, i5 );
nand ( wi9, i2, i7 );
nor ( wi10, i9, i11 );
or ( wi11, i4, i5 );
xor ( wi12, i10, i15 );
and ( wi13, i13, i17 );
xor ( wi14, i11, i18 );
or ( wi15, i0, i12 );
or ( wi16, i1, i4 );
and ( wi17, i12, i18 );
or ( wi18, i1, i6 );
or ( wi19, i13, i14 );
and ( wi20, i1, i17 );
or ( wi21, i0, i3 );
nor ( wi22, i1, i15 );
nor ( wi23, wi1, wi12 );
nor ( wi24, wi1, wi17 );
nor ( wi25, wi0, wi20 );
xor ( wi26, wi1, wi4 );
xor ( wi27, wi20, wi21 );
nand ( wi28, wi14, wi15 );
nand ( wi29, wi3, wi12 );
nor ( wi30, wi5, wi17 );
xor ( wi31, wi5, wi10 );
or ( wi32, wi13, wi18 );
or ( wi33, wi0, wi9 );
or ( wi34, wi5, wi13 );
or ( wi35, wi5, wi21 );
xor ( wi36, wi15, wi17 );
and ( wi37, wi1, wi4 );
nand ( wi38, wi29, wi30 );
nor ( wi39, wi11, wi25 );
nor ( wi40, wi11, wi32 );
xor ( wi41, wi19, wi31 );
nor ( wi42, wi6, wi11 );
or ( wi43, wi5, wi9 );
or ( wi44, wi7, wi28 );
and ( wi45, wi13, wi17 );
and ( wi46, wi5, wi18 );
nand ( wi47, wi4, wi14 );
or ( wi48, wi6, wi16 );
and ( wi49, wi17, wi22 );
and ( wi50, wi7, wi11 );
xor ( wi51, wi1, wi17 );
or ( wi52, wi20, wi21 );
nand ( wi53, wi27, wi28 );
and ( wi54, wi7, wi12 );
nor ( wi55, wi5, wi28 );
xor ( wi56, wi0, wi13 );
nor ( wi57, wi2, wi18 );
xor ( wi58, wi0, wi5 );
or ( wi59, wi18, wi23 );
nand ( wi60, wi29, wi42 );
and ( wi61, wi16, wi56 );
and ( wi62, wi29, wi45 );
xor ( wi63, wi18, wi40 );
or ( wi64, wi6, wi40 );
xor ( wi65, wi32, wi35 );
and ( wi66, wi30, wi37 );
nand ( wi67, wi31, wi46 );
xor ( wi68, wi34, wi56 );
nor ( wi69, wi8, wi20 );
and ( wi70, wi3, wi11 );
or ( wi71, wi22, wi57 );
nor ( wi72, wi55, wi56 );
or ( wi73, wi5, wi56 );
and ( wi74, wi32, wi57 );
nand ( wi75, wi2, wi55 );
or ( wi76, wi7, wi23 );
and ( wi77, wi29, wi56 );
or ( wi78, wi26, wi49 );
and ( wi79, wi31, wi35 );
or ( wi80, wi7, wi54 );
and ( wi81, wi39, wi44 );
or ( wi82, wi25, wi34 );
or ( wi83, wi11, wi23 );
nor ( wi84, wi10, wi17 );
nand ( wi85, wi10, wi11 );
or ( wi86, wi40, wi41 );
or ( wi87, wi8, wi56 );
xor ( wi88, wi24, wi54 );
xor ( wi89, wi32, wi47 );
or ( wi90, wi24, wi48 );
nand ( wi91, wi26, wi52 );
and ( wi92, wi43, wi44 );
xor ( wi93, wi22, wi40 );
nand ( wi94, wi18, wi47 );
and ( wi95, wi17, wi18 );
nand ( wi96, wi38, wi48 );
or ( wi97, wi27, wi57 );
nand ( wi98, wi18, wi34 );
and ( wi99, wi28, wi56 );
nor ( wi100, wi4, wi57 );
and ( wi101, wi15, wi54 );
and ( wi102, wi19, wi27 );
nor ( wi103, wi27, wi33 );
xor ( wi104, wi1, wi48 );
and ( wi105, wi39, wi40 );
nand ( wi106, wi9, wi45 );
xor ( wi107, wi1, wi45 );
nand ( wi108, wi14, wi16 );
xor ( wi109, wi30, wi51 );
nand ( wi110, wi27, wi31 );
nand ( wi111, wi3, wi50 );
nand ( wi112, wi51, wi55 );
and ( wi113, wi10, wi45 );
xor ( wi114, wi21, wi39 );
xor ( wi115, wi7, wi50 );
xor ( wi116, wi1, wi2 );
or ( wi117, wi29, wi49 );
xor ( wi118, wi16, wi58 );
and ( wi119, wi17, wi47 );
and ( wi120, wi35, wi45 );
and ( wi121, wi24, wi28 );
xor ( wi122, wi23, wi29 );
nor ( wi123, wi6, wi36 );
xor ( wi124, wi23, wi54 );
and ( wi125, wi11, wi30 );
or ( wi126, wi10, wi19 );
and ( wi127, wi17, wi26 );
xor ( wi128, wi17, wi30 );
and ( wi129, wi26, wi45 );
xor ( wi130, wi11, wi36 );
and ( wi131, wi3, wi26 );
or ( wi132, wi31, wi57 );
nor ( wi133, wi24, wi56 );
or ( wi134, wi15, wi40 );
xor ( wi135, wi56, wi58 );
nand ( wi136, wi9, wi54 );
nand ( wi137, wi27, wi51 );
or ( wi138, wi5, wi41 );
and ( wi139, wi1, wi13 );
nand ( wi140, wi6, wi50 );
nor ( wi141, wi0, wi5 );
and ( wi142, wi27, wi54 );
nand ( wi143, wi40, wi47 );
and ( wi144, wi28, wi42 );
or ( wi145, wi48, wi115 );
and ( wi146, wi101, wi143 );
nor ( wi147, wi8, wi33 );
nand ( wi148, wi43, wi133 );
or ( wi149, wi77, wi103 );
or ( wi150, wi12, wi46 );
and ( wi151, wi65, wi85 );
xor ( wi152, wi128, wi129 );
nor ( wi153, wi47, wi57 );
nand ( wi154, wi123, wi124 );
nand ( wi155, wi48, wi136 );
or ( wi156, wi4, wi59 );
xor ( wi157, wi51, wi99 );
or ( wi158, wi10, wi129 );
or ( wi159, wi19, wi115 );
or ( wi160, wi60, wi126 );
nor ( wi161, wi24, wi140 );
xor ( wi162, wi6, wi20 );
nor ( wi163, wi33, wi124 );
and ( wi164, wi26, wi135 );
or ( wi165, wi75, wi130 );
nand ( wi166, wi10, wi50 );
and ( wi167, wi16, wi43 );
or ( wi168, wi54, wi115 );
nand ( wi169, wi27, wi139 );
nand ( wi170, wi64, wi129 );
and ( wi171, wi33, wi74 );
and ( wi172, wi71, wi120 );
nand ( wi173, wi106, wi110 );
xor ( wi174, wi6, wi38 );
nand ( wi175, wi47, wi94 );
xor ( wi176, wi97, wi135 );
nand ( wi177, wi100, wi117 );
nand ( wi178, wi42, wi110 );
and ( wi179, wi40, wi58 );
and ( wi180, wi16, wi29 );
or ( wi181, wi36, wi67 );
and ( wi182, wi24, wi126 );
or ( wi183, wi22, wi80 );
and ( wi184, wi13, wi44 );
nand ( wi185, wi0, wi108 );
and ( wi186, wi104, wi114 );
and ( wi187, wi113, wi134 );
xor ( wi188, wi20, wi36 );
nor ( wi189, wi100, wi125 );
or ( wi190, wi21, wi23 );
nand ( wi191, wi64, wi67 );
or ( wi192, wi3, wi43 );
or ( wi193, wi21, wi56 );
nor ( wi194, wi24, wi64 );
xor ( wi195, wi10, wi128 );
nor ( wi196, wi98, wi141 );
xor ( wi197, wi78, wi119 );
xor ( wi198, wi63, wi67 );
or ( wi199, wi94, wi104 );
or ( wi200, wi22, wi35 );
xor ( wi201, wi82, wi106 );
xor ( wi202, wi20, wi86 );
xor ( wi203, wi14, wi76 );
nor ( wi204, wi8, wi26 );
nand ( wi205, wi67, wi69 );
nor ( wi206, wi88, wi140 );
xor ( wi207, wi40, wi143 );
nor ( wi208, wi14, wi25 );
or ( wi209, wi37, wi91 );
and ( wi210, wi47, wi117 );
xor ( wi211, wi40, wi69 );
or ( wi212, wi105, wi111 );
and ( wi213, wi97, wi107 );
nor ( wi214, wi35, wi81 );
nand ( wi215, wi82, wi86 );
xor ( wi216, wi36, wi143 );
xor ( wi217, wi17, wi102 );
and ( wi218, wi123, wi127 );
or ( wi219, wi30, wi31 );
or ( wi220, wi46, wi89 );
and ( wi221, wi44, wi75 );
nand ( wi222, wi103, wi131 );
or ( wi223, wi16, wi30 );
nand ( wi224, wi17, wi52 );
or ( wi225, wi82, wi116 );
xor ( wi226, wi38, wi85 );
xor ( wi227, wi62, wi142 );
or ( wi228, wi119, wi120 );
or ( wi229, wi68, wi113 );
nor ( wi230, wi97, wi112 );
and ( wi231, wi5, wi89 );
xor ( wi232, wi16, wi39 );
and ( wi233, wi101, wi122 );
nand ( wi234, wi94, wi110 );
xor ( wi235, wi50, wi79 );
or ( wi236, wi90, wi139 );
or ( wi237, wi68, wi95 );
or ( wi238, wi20, wi120 );
or ( wi239, wi14, wi88 );
nor ( wi240, wi81, wi98 );
or ( wi241, wi39, wi77 );
or ( wi242, wi45, wi112 );
or ( wi243, wi116, wi136 );
nor ( wi244, wi62, wi105 );
or ( wi245, wi5, wi108 );
nand ( wi246, wi5, wi93 );
nand ( wi247, wi1, wi10 );
nor ( wi248, wi83, wi143 );
nand ( wi249, wi22, wi118 );
xor ( wi250, wi1, wi78 );
and ( wi251, wi66, wi82 );
and ( wi252, wi3, wi54 );
and ( wi253, wi26, wi57 );
and ( wi254, wi107, wi125 );
xor ( wi255, wi19, wi141 );
xor ( wi256, wi58, wi116 );
or ( wi257, wi7, wi136 );
nand ( wi258, wi26, wi105 );
or ( wi259, wi23, wi89 );
nand ( wi260, wi84, wi138 );
nand ( wi261, wi109, wi111 );
and ( wi262, wi1, wi116 );
xor ( wi263, wi63, wi64 );
or ( wi264, wi27, wi59 );
or ( wi265, wi53, wi91 );
nor ( wi266, wi108, wi139 );
xor ( wi267, wi29, wi31 );
nand ( wi268, wi133, wi139 );
nor ( wi269, wi8, wi13 );
nor ( wi270, wi8, wi46 );
nor ( wi271, wi78, wi121 );
xor ( wi272, wi56, wi57 );
or ( wi273, wi57, wi118 );
nand ( wi274, wi47, wi112 );
nor ( wi275, wi6, wi108 );
or ( wi276, wi14, wi39 );
xor ( wi277, wi31, wi40 );
and ( wi278, wi6, wi23 );
or ( wi279, wi84, wi121 );
or ( wi280, wi24, wi52 );
xor ( wi281, wi20, wi113 );
and ( wi282, wi54, wi132 );
xor ( wi283, wi18, wi66 );
and ( wi284, wi110, wi116 );
or ( wi285, wi1, wi94 );
nor ( wi286, wi86, wi134 );
or ( wi287, wi79, wi142 );
nor ( wi288, wi120, wi123 );
and ( wi289, wi125, wi140 );
and ( wi290, wi38, wi117 );
nand ( wi291, wi29, wi100 );
nor ( wi292, wi62, wi90 );
or ( wi293, wi46, wi116 );
nand ( wi294, wi20, wi99 );
and ( wi295, wi60, wi79 );
xor ( wi296, wi3, wi39 );
xor ( wi297, wi115, wi132 );
nor ( wi298, wi50, wi142 );
nand ( wi299, wi2, wi103 );
xor ( wi300, wi99, wi108 );
nor ( wi301, wi4, wi31 );
nor ( wi302, wi35, wi112 );
nor ( wi303, wi18, wi53 );
nand ( wi304, wi50, wi116 );
and ( wi305, wi77, wi135 );
or ( wi306, wi31, wi51 );
nor ( wi307, wi26, wi58 );
and ( wi308, wi129, wi138 );
nand ( wi309, wi31, wi85 );
and ( wi310, wi113, wi120 );
nor ( wi311, wi33, wi112 );
or ( wi312, wi121, wi129 );
nand ( wi313, wi38, wi59 );
nor ( wi314, wi59, wi125 );
and ( wi315, wi62, wi83 );
xor ( wi316, wi119, wi135 );
and ( wi317, wi115, wi130 );
nor ( wi318, wi57, wi129 );
xor ( wi319, wi106, wi131 );
or ( wi320, wi86, wi109 );
nor ( wi321, wi5, wi30 );
or ( wi322, wi32, wi133 );
nor ( wi323, wi71, wi79 );
nand ( wi324, wi67, wi110 );
nor ( wi325, wi128, wi140 );
nand ( wi326, wi54, wi104 );
nand ( wi327, wi37, wi116 );
xor ( wi328, wi66, wi71 );
or ( wi329, wi9, wi110 );
or ( wi330, wi43, wi70 );
or ( wi331, wi48, wi84 );
or ( wi332, wi18, wi86 );
and ( wi333, wi46, wi90 );
xor ( wi334, wi40, wi141 );
or ( wi335, wi67, wi74 );
and ( wi336, wi28, wi35 );
or ( wi337, wi93, wi112 );
or ( wi338, wi23, wi63 );
xor ( wi339, wi133, wi134 );
and ( wi340, wi25, wi78 );
and ( wi341, wi43, wi118 );
xor ( wi342, wi56, wi114 );
or ( wi343, wi50, wi69 );
or ( wi344, wi74, wi141 );
nand ( wi345, wi30, wi103 );
and ( wi346, wi79, wi135 );
nand ( wi347, wi41, wi90 );
xor ( wi348, wi137, wi141 );
and ( wi349, wi65, wi118 );
xor ( wi350, wi36, wi100 );
nor ( wi351, wi81, wi100 );
xor ( wi352, wi45, wi57 );
nor ( wi353, wi9, wi89 );
xor ( wi354, wi22, wi46 );
xor ( wi355, wi112, wi143 );
and ( wi356, wi34, wi128 );
nand ( wi357, wi14, wi32 );
nand ( wi358, wi29, wi112 );
nor ( wi359, wi5, wi134 );
or ( wi360, wi69, wi89 );
nor ( wi361, wi87, wi108 );
or ( wi362, wi19, wi88 );
nand ( wi363, wi37, wi82 );
nor ( wi364, wi5, wi106 );
nand ( wi365, wi0, wi97 );
and ( wi366, wi69, wi108 );
nor ( wi367, wi34, wi110 );
xor ( wi368, wi13, wi19 );
nand ( wi369, wi25, wi119 );
and ( wi370, wi92, wi137 );
xor ( wi371, wi88, wi126 );
xor ( wi372, wi40, wi82 );
xor ( wi373, wi19, wi109 );
xor ( wi374, wi52, wi142 );
nor ( wi375, wi5, wi64 );
and ( wi376, wi112, wi120 );
nand ( wi377, wi30, wi69 );
and ( wi378, wi5, wi69 );
and ( wi379, wi55, wi133 );
and ( wi380, wi15, wi73 );
nor ( wi381, wi10, wi117 );
nor ( wi382, wi30, wi65 );
or ( wi383, wi21, wi46 );
or ( wi384, wi103, wi141 );
and ( wi385, wi56, wi122 );
nand ( wi386, wi73, wi109 );
nor ( wi387, wi28, wi111 );
nand ( wi388, wi40, wi110 );
and ( wi389, wi84, wi92 );
xor ( wi390, wi6, wi75 );
xor ( wi391, wi40, wi111 );
nand ( wi392, wi99, wi118 );
nand ( wi393, wi1, wi126 );
xor ( wi394, wi0, wi79 );
or ( wi395, wi62, wi100 );
and ( wi396, wi99, wi121 );
nor ( wi397, wi19, wi130 );
and ( wi398, wi9, wi95 );
nand ( wi399, wi8, wi82 );
nand ( wi400, wi36, wi140 );
or ( wi401, wi92, wi118 );
nand ( wi402, wi33, wi107 );
nand ( wi403, wi23, wi135 );
nor ( wi404, wi52, wi95 );
xor ( wi405, wi14, wi48 );
and ( wi406, wi36, wi75 );
nand ( wi407, wi37, wi90 );
and ( wi408, wi32, wi113 );
nor ( wi409, wi118, wi127 );
nand ( wi410, wi48, wi109 );
nor ( wi411, wi39, wi139 );
or ( wi412, wi11, wi12 );
xor ( wi413, wi0, wi87 );
nor ( wi414, wi3, wi124 );
or ( wi415, wi3, wi126 );
nand ( wi416, wi21, wi44 );
nor ( wi417, wi13, wi56 );
xor ( wi418, wi52, wi89 );
and ( wi419, wi65, wi67 );
or ( wi420, wi6, wi64 );
or ( wi421, wi60, wi107 );
nor ( wi422, wi112, wi129 );
and ( wi423, wi35, wi132 );
nor ( wi424, wi51, wi140 );
xor ( wi425, wi93, wi108 );
nor ( wi426, wi2, wi139 );
nand ( wi427, wi89, wi113 );
nand ( wi428, wi40, wi102 );
nor ( wi429, wi13, wi53 );
or ( wi430, wi26, wi63 );
and ( wi431, wi106, wi136 );
nor ( wi432, wi45, wi125 );
nand ( wi433, wi56, wi58 );
xor ( wi434, wi15, wi134 );
xor ( wi435, wi5, wi83 );
xor ( wi436, wi57, wi84 );
and ( wi437, wi13, wi120 );
nand ( wi438, wi5, wi97 );
or ( wi439, wi38, wi56 );
xor ( wi440, wi11, wi20 );
and ( wi441, wi13, wi101 );
nor ( wi442, wi30, wi102 );
xor ( wi443, wi56, wi101 );
xor ( wi444, wi98, wi129 );
xor ( wi445, wi8, wi68 );
and ( wi446, wi115, wi126 );
nor ( wi447, wi81, wi143 );
and ( wi448, wi93, wi104 );
or ( wi449, wi17, wi83 );
and ( wi450, wi99, wi120 );
or ( wi451, wi55, wi111 );
nor ( wi452, wi38, wi86 );
nor ( wi453, wi44, wi130 );
xor ( wi454, wi105, wi107 );
or ( wi455, wi30, wi143 );
nand ( wi456, wi89, wi136 );
or ( wi457, wi116, wi131 );
nor ( wi458, wi60, wi116 );
and ( wi459, wi137, wi143 );
nand ( wi460, wi0, wi103 );
and ( wi461, wi126, wi140 );
nand ( wi462, wi23, wi99 );
nand ( wi463, wi85, wi130 );
and ( wi464, wi7, wi73 );
or ( wi465, wi27, wi44 );
nand ( wi466, wi12, wi75 );
and ( wi467, wi5, wi43 );
nor ( wi468, wi112, wi141 );
and ( wi469, wi39, wi114 );
nand ( wi470, wi4, wi99 );
or ( wi471, wi29, wi136 );
nand ( wi472, wi55, wi106 );
nand ( wi473, wi8, wi63 );
xor ( wi474, wi5, wi122 );
and ( wi475, wi18, wi102 );
and ( wi476, wi40, wi108 );
nand ( wi477, wi30, wi86 );
nor ( wi478, wi83, wi141 );
nand ( wi479, wi133, wi143 );
or ( wi480, wi21, wi67 );
xor ( wi481, wi6, wi116 );
or ( wi482, wi65, wi117 );
and ( wi483, wi81, wi122 );
or ( wi484, wi4, wi85 );
nand ( wi485, wi21, wi93 );
nor ( wi486, wi37, wi76 );
nand ( wi487, wi52, wi96 );
xor ( wi488, wi70, wi101 );
and ( wi489, wi121, wi134 );
nand ( wi490, wi7, wi54 );
or ( wi491, wi81, wi115 );
or ( wi492, wi7, wi9 );
or ( wi493, wi47, wi130 );
nor ( wi494, wi25, wi132 );
xor ( wi495, wi60, wi80 );
or ( wi496, wi106, wi121 );
and ( wi497, wi23, wi138 );
nand ( wi498, wi43, wi121 );
or ( wi499, wi8, wi69 );
and ( wi500, wi64, wi120 );
or ( wi501, wi60, wi113 );
nor ( wi502, wi18, wi40 );
and ( wi503, wi5, wi139 );
nor ( wi504, wi20, wi69 );
and ( wi505, wi48, wi60 );
nor ( wi506, wi44, wi98 );
or ( wi507, wi29, wi76 );
nor ( wi508, wi116, wi142 );
nand ( wi509, wi46, wi91 );
nor ( wi510, wi48, wi127 );
and ( wi511, wi7, wi21 );
and ( wi512, wi72, wi82 );
or ( wi513, wi91, wi112 );
or ( wi514, wi111, wi117 );
nor ( wi515, wi123, wi139 );
or ( wi516, wi88, wi130 );
xor ( wi517, wi62, wi123 );
or ( wi518, wi19, wi120 );
and ( wi519, wi61, wi66 );
xor ( wi520, wi44, wi133 );
nand ( wi521, wi102, wi129 );
nor ( wi522, wi7, wi14 );
and ( wi523, wi43, wi80 );
or ( wi524, wi62, wi124 );
or ( wi525, wi26, wi97 );
nor ( wi526, wi33, wi62 );
nor ( wi527, wi90, wi118 );
nor ( wi528, wi82, wi89 );
and ( wi529, wi14, wi50 );
xor ( wi530, wi26, wi53 );
xor ( wi531, wi40, wi113 );
xor ( wi532, wi17, wi99 );
nor ( wi533, wi12, wi130 );
nand ( wi534, wi25, wi73 );
and ( wi535, wi73, wi76 );
nor ( wi536, wi19, wi110 );
nor ( wi537, wi60, wi102 );
or ( wi538, wi31, wi53 );
nand ( wi539, wi112, wi140 );
nand ( wi540, wi50, wi114 );
nor ( wi541, wi27, wi38 );
nor ( wi542, wi55, wi93 );
nand ( wi543, wi31, wi99 );
and ( wi544, wi32, wi34 );
nor ( wi545, wi48, wi140 );
xor ( wi546, wi59, wi141 );
xor ( wi547, wi1, wi109 );
and ( wi548, wi10, wi48 );
nand ( wi549, wi21, wi28 );
or ( wi550, wi64, wi143 );
nand ( wi551, wi1, wi8 );
nand ( wi552, wi110, wi114 );
or ( wi553, wi98, wi101 );
and ( wi554, wi40, wi128 );
xor ( wi555, wi17, wi139 );
nor ( wi556, wi59, wi126 );
nand ( wi557, wi22, wi98 );
or ( wi558, wi45, wi91 );
nand ( wi559, wi16, wi58 );
nor ( wi560, wi30, wi131 );
nand ( wi561, wi109, wi134 );
or ( wi562, wi76, wi79 );
nand ( wi563, wi49, wi124 );
and ( wi564, wi8, wi94 );
xor ( wi565, wi37, wi107 );
or ( wi566, wi53, wi74 );
nor ( wi567, wi27, wi142 );
or ( wi568, wi84, wi114 );
or ( wi569, wi87, wi132 );
or ( wi570, wi99, wi122 );
and ( wi571, wi103, wi134 );
or ( wi572, wi5, wi95 );
nor ( wi573, wi16, wi86 );
nor ( wi574, wi78, wi97 );
xor ( wi575, wi14, wi118 );
and ( wi576, wi10, wi45 );
or ( wi577, wi70, wi89 );
nand ( wi578, wi110, wi142 );
nand ( wi579, wi43, wi47 );
xor ( wi580, wi3, wi4 );
xor ( wi581, wi96, wi139 );
nor ( wi582, wi10, wi125 );
xor ( wi583, wi28, wi115 );
nand ( wi584, wi21, wi70 );
or ( wi585, wi98, wi137 );
and ( wi586, wi39, wi63 );
and ( wi587, wi51, wi101 );
xor ( wi588, wi57, wi98 );
nor ( wi589, wi58, wi115 );
or ( wi590, wi46, wi142 );
xor ( wi591, wi15, wi27 );
nor ( wi592, wi13, wi33 );
nor ( wi593, wi65, wi90 );
or ( wi594, wi31, wi143 );
nor ( wi595, wi56, wi83 );
nand ( wi596, wi21, wi103 );
nand ( wi597, wi82, wi136 );
xor ( wi598, wi64, wi86 );
nand ( wi599, wi36, wi87 );
nor ( wi600, wi2, wi19 );
nor ( wi601, wi63, wi78 );
or ( wi602, wi89, wi123 );
or ( wi603, wi24, wi49 );
or ( wi604, wi31, wi80 );
nand ( wi605, wi33, wi58 );
and ( wi606, wi0, wi138 );
or ( wi607, wi111, wi123 );
or ( wi608, wi21, wi54 );
nor ( wi609, wi114, wi119 );
nand ( wi610, wi34, wi44 );
nand ( wi611, wi64, wi141 );
and ( wi612, wi29, wi138 );
nor ( wi613, wi13, wi140 );
xor ( wi614, wi2, wi73 );
nand ( wi615, wi68, wi130 );
or ( wi616, wi14, wi104 );
or ( wi617, wi5, wi67 );
nand ( wi618, wi54, wi122 );
nor ( wi619, wi1, wi114 );
nand ( wi620, wi4, wi122 );
nand ( wi621, wi14, wi138 );
or ( wi622, wi97, wi142 );
nand ( wi623, wi40, wi50 );
or ( wi624, wi64, wi90 );
or ( wi625, wi91, wi136 );
and ( wi626, wi38, wi141 );
nand ( wi627, wi52, wi58 );
and ( wi628, wi30, wi122 );
nor ( wi629, wi31, wi105 );
nand ( wi630, wi63, wi101 );
nand ( wi631, wi93, wi115 );
and ( wi632, wi65, wi140 );
nand ( wi633, wi65, wi120 );
nand ( wi634, wi59, wi90 );
or ( wi635, wi15, wi123 );
nand ( wi636, wi40, wi59 );
nor ( wi637, wi42, wi77 );
nand ( wi638, wi36, wi54 );
and ( wi639, wi72, wi88 );
and ( wi640, wi47, wi68 );
nor ( wi641, wi120, wi141 );
nor ( wi642, wi15, wi51 );
and ( wi643, wi13, wi74 );
nor ( wi644, wi7, wi72 );
nand ( wi645, wi42, wi62 );
xor ( wi646, wi49, wi68 );
xor ( wi647, wi96, wi140 );
nor ( wi648, wi0, wi21 );
and ( wi649, wi101, wi109 );
and ( wi650, wi42, wi79 );
nor ( wi651, wi45, wi129 );
nor ( wi652, wi80, wi84 );
nand ( wi653, wi52, wi126 );
or ( wi654, wi26, wi99 );
nor ( wi655, wi15, wi119 );
nand ( wi656, wi3, wi97 );
nor ( wi657, wi34, wi61 );
xor ( wi658, wi81, wi114 );
nor ( ou0, i1, i0 );
nor ( ou1, i3, i16 );
xor ( ou2, i9, i17 );
nand ( ou3, i0, i7 );
or ( ou4, i13, i16 );
nor ( ou5, i1, i0 );
or ( ou6, i3, i11 );
and ( ou7, i5, i10 );
nor ( ou8, i11, i7 );
or ( ou9, i15, i18 );
nor ( ou10, i9, i17 );

endmodule
